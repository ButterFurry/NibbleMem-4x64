* NGSPICE file created from nibble_mem.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR Q CLK R S D gnd vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

.subckt nibble_mem vdd gnd clk rst_n din[0] din[1] din[2] din[3] store next prev dout[0]
+ dout[1] dout[2] dout[3] addr[0] addr[1] addr[2] addr[3] addr[4] addr[5]
XFILL_65_DFFSR_227 gnd vdd FILL
XFILL_87_DFFSR_69 gnd vdd FILL
XFILL_16_DFFSR_25 gnd vdd FILL
XFILL_9_6_0 gnd vdd FILL
XFILL_16_DFFSR_36 gnd vdd FILL
XFILL_65_DFFSR_238 gnd vdd FILL
XFILL_65_DFFSR_249 gnd vdd FILL
XFILL_19_NOR3X1_15 gnd vdd FILL
XFILL_16_DFFSR_47 gnd vdd FILL
XFILL_16_DFFSR_58 gnd vdd FILL
XFILL_19_NOR3X1_26 gnd vdd FILL
XFILL_16_DFFSR_69 gnd vdd FILL
XFILL_19_NOR3X1_37 gnd vdd FILL
XFILL_19_NOR3X1_48 gnd vdd FILL
XFILL_69_DFFSR_204 gnd vdd FILL
XFILL_56_DFFSR_13 gnd vdd FILL
XFILL_69_DFFSR_215 gnd vdd FILL
XFILL_13_CLKBUF1_40 gnd vdd FILL
XFILL_56_DFFSR_24 gnd vdd FILL
XFILL_69_DFFSR_226 gnd vdd FILL
XFILL_56_DFFSR_35 gnd vdd FILL
XFILL_48_1_2 gnd vdd FILL
XFILL_69_DFFSR_237 gnd vdd FILL
XFILL_56_DFFSR_46 gnd vdd FILL
XFILL_69_DFFSR_248 gnd vdd FILL
XFILL_69_DFFSR_259 gnd vdd FILL
XFILL_56_DFFSR_57 gnd vdd FILL
XFILL_56_DFFSR_68 gnd vdd FILL
XFILL_56_DFFSR_79 gnd vdd FILL
XFILL_17_5_0 gnd vdd FILL
XFILL_54_DFFSR_6 gnd vdd FILL
XFILL_25_DFFSR_12 gnd vdd FILL
XFILL_25_DFFSR_23 gnd vdd FILL
XFILL_25_DFFSR_34 gnd vdd FILL
XFILL_25_DFFSR_45 gnd vdd FILL
XFILL_25_DFFSR_56 gnd vdd FILL
XFILL_11_NOR2X1_180 gnd vdd FILL
XFILL_25_DFFSR_67 gnd vdd FILL
XFILL_11_NOR2X1_191 gnd vdd FILL
XFILL_25_DFFSR_78 gnd vdd FILL
XFILL_31_0_2 gnd vdd FILL
XFILL_25_DFFSR_89 gnd vdd FILL
XFILL_65_DFFSR_11 gnd vdd FILL
XFILL_65_DFFSR_22 gnd vdd FILL
XFILL_50_DFFSR_260 gnd vdd FILL
XFILL_50_DFFSR_271 gnd vdd FILL
XFILL_65_DFFSR_33 gnd vdd FILL
XFILL_65_DFFSR_44 gnd vdd FILL
XFILL_0_MUX2X1_9 gnd vdd FILL
XFILL_65_DFFSR_55 gnd vdd FILL
XFILL_65_DFFSR_66 gnd vdd FILL
XFILL_65_DFFSR_77 gnd vdd FILL
XFILL_65_DFFSR_88 gnd vdd FILL
XFILL_65_DFFSR_99 gnd vdd FILL
XFILL_15_NAND3X1_107 gnd vdd FILL
XFILL_15_NAND3X1_118 gnd vdd FILL
XFILL_8_DFFSR_13 gnd vdd FILL
XFILL_54_DFFSR_270 gnd vdd FILL
XFILL_15_NAND3X1_129 gnd vdd FILL
XFILL_8_DFFSR_24 gnd vdd FILL
XFILL_19_DFFSR_9 gnd vdd FILL
XFILL_8_DFFSR_35 gnd vdd FILL
XFILL_34_DFFSR_10 gnd vdd FILL
XFILL_34_DFFSR_21 gnd vdd FILL
XFILL_8_DFFSR_46 gnd vdd FILL
XFILL_11_MUX2X1_120 gnd vdd FILL
XFILL_8_DFFSR_57 gnd vdd FILL
XFILL_34_DFFSR_32 gnd vdd FILL
XFILL_11_MUX2X1_131 gnd vdd FILL
XFILL_34_DFFSR_43 gnd vdd FILL
XFILL_8_DFFSR_68 gnd vdd FILL
XFILL_8_DFFSR_79 gnd vdd FILL
XFILL_11_MUX2X1_142 gnd vdd FILL
XFILL_34_DFFSR_54 gnd vdd FILL
XFILL_11_MUX2X1_153 gnd vdd FILL
XFILL_34_DFFSR_65 gnd vdd FILL
XFILL_34_DFFSR_76 gnd vdd FILL
XFILL_81_DFFSR_170 gnd vdd FILL
XFILL_11_MUX2X1_164 gnd vdd FILL
XFILL_11_MUX2X1_175 gnd vdd FILL
XFILL_81_DFFSR_181 gnd vdd FILL
XFILL_11_MUX2X1_186 gnd vdd FILL
XFILL_34_DFFSR_87 gnd vdd FILL
XFILL_34_DFFSR_98 gnd vdd FILL
XFILL_81_DFFSR_192 gnd vdd FILL
XFILL_32_DFFSR_205 gnd vdd FILL
XFILL_74_DFFSR_20 gnd vdd FILL
XFILL_32_DFFSR_216 gnd vdd FILL
XFILL_74_DFFSR_31 gnd vdd FILL
XFILL_32_DFFSR_227 gnd vdd FILL
XFILL_1_DFFSR_240 gnd vdd FILL
XFILL_1_DFFSR_251 gnd vdd FILL
XFILL_32_DFFSR_238 gnd vdd FILL
XFILL_74_DFFSR_42 gnd vdd FILL
XFILL_32_DFFSR_249 gnd vdd FILL
XFILL_74_DFFSR_53 gnd vdd FILL
XFILL_1_DFFSR_262 gnd vdd FILL
XFILL_74_DFFSR_64 gnd vdd FILL
XFILL_1_DFFSR_273 gnd vdd FILL
XFILL_74_DFFSR_75 gnd vdd FILL
XFILL_85_DFFSR_180 gnd vdd FILL
XFILL_74_DFFSR_86 gnd vdd FILL
XFILL_39_1_2 gnd vdd FILL
XFILL_85_DFFSR_191 gnd vdd FILL
XFILL_36_DFFSR_204 gnd vdd FILL
XFILL_74_DFFSR_97 gnd vdd FILL
XFILL_36_DFFSR_215 gnd vdd FILL
XFILL_36_DFFSR_226 gnd vdd FILL
XFILL_36_DFFSR_237 gnd vdd FILL
XFILL_5_DFFSR_250 gnd vdd FILL
XFILL_36_DFFSR_248 gnd vdd FILL
XFILL_5_DFFSR_261 gnd vdd FILL
XFILL_5_DFFSR_272 gnd vdd FILL
XFILL_43_DFFSR_30 gnd vdd FILL
XFILL_36_DFFSR_259 gnd vdd FILL
XFILL_43_DFFSR_41 gnd vdd FILL
XFILL_2_MUX2X1_17 gnd vdd FILL
XFILL_14_NOR3X1_5 gnd vdd FILL
XFILL_2_MUX2X1_28 gnd vdd FILL
XFILL_63_DFFSR_104 gnd vdd FILL
XFILL_43_DFFSR_52 gnd vdd FILL
XFILL_43_DFFSR_63 gnd vdd FILL
XFILL_2_MUX2X1_39 gnd vdd FILL
XFILL_63_DFFSR_115 gnd vdd FILL
XFILL_43_DFFSR_74 gnd vdd FILL
XFILL_63_DFFSR_126 gnd vdd FILL
XFILL_43_DFFSR_85 gnd vdd FILL
XFILL_63_DFFSR_137 gnd vdd FILL
XFILL_43_DFFSR_96 gnd vdd FILL
XFILL_63_DFFSR_148 gnd vdd FILL
XFILL_10_NAND3X1_103 gnd vdd FILL
XFILL_9_DFFSR_260 gnd vdd FILL
XFILL_10_NAND3X1_114 gnd vdd FILL
XFILL_63_DFFSR_159 gnd vdd FILL
XFILL_9_DFFSR_271 gnd vdd FILL
XFILL_10_NAND3X1_125 gnd vdd FILL
XFILL_83_DFFSR_40 gnd vdd FILL
XFILL_50_3_0 gnd vdd FILL
XFILL_6_MUX2X1_16 gnd vdd FILL
XFILL_83_DFFSR_51 gnd vdd FILL
XFILL_6_MUX2X1_27 gnd vdd FILL
XFILL_67_DFFSR_103 gnd vdd FILL
XFILL_22_0_2 gnd vdd FILL
XFILL_6_MUX2X1_38 gnd vdd FILL
XFILL_67_DFFSR_114 gnd vdd FILL
XFILL_83_DFFSR_62 gnd vdd FILL
XFILL_83_DFFSR_73 gnd vdd FILL
XFILL_6_MUX2X1_49 gnd vdd FILL
XFILL_67_DFFSR_125 gnd vdd FILL
XFILL_67_DFFSR_136 gnd vdd FILL
XFILL_83_DFFSR_84 gnd vdd FILL
XFILL_12_DFFSR_40 gnd vdd FILL
XFILL_83_DFFSR_95 gnd vdd FILL
XFILL_12_DFFSR_51 gnd vdd FILL
XFILL_10_OAI21X1_4 gnd vdd FILL
XFILL_14_NAND3X1_12 gnd vdd FILL
XFILL_67_DFFSR_147 gnd vdd FILL
XFILL_67_DFFSR_158 gnd vdd FILL
XFILL_1_MUX2X1_170 gnd vdd FILL
XFILL_14_NAND3X1_23 gnd vdd FILL
XFILL_12_DFFSR_62 gnd vdd FILL
XFILL_12_DFFSR_73 gnd vdd FILL
XFILL_67_DFFSR_169 gnd vdd FILL
XFILL_14_NAND3X1_34 gnd vdd FILL
XFILL_1_MUX2X1_181 gnd vdd FILL
XFILL_12_DFFSR_84 gnd vdd FILL
XFILL_13_BUFX4_9 gnd vdd FILL
XFILL_14_NAND3X1_45 gnd vdd FILL
XFILL_1_MUX2X1_192 gnd vdd FILL
XFILL_12_DFFSR_95 gnd vdd FILL
XFILL_14_NAND3X1_56 gnd vdd FILL
XFILL_34_CLKBUF1_12 gnd vdd FILL
XFILL_14_NAND3X1_67 gnd vdd FILL
XFILL_34_CLKBUF1_23 gnd vdd FILL
XFILL_14_NAND3X1_78 gnd vdd FILL
XFILL_34_CLKBUF1_34 gnd vdd FILL
XFILL_23_NOR3X1_3 gnd vdd FILL
XFILL_14_NAND3X1_89 gnd vdd FILL
XFILL_52_DFFSR_50 gnd vdd FILL
XFILL_14_OAI21X1_3 gnd vdd FILL
XFILL_1_NAND3X1_108 gnd vdd FILL
XFILL_52_DFFSR_61 gnd vdd FILL
XFILL_1_NAND3X1_119 gnd vdd FILL
XFILL_11_NOR2X1_50 gnd vdd FILL
XFILL_52_DFFSR_72 gnd vdd FILL
XFILL_52_DFFSR_83 gnd vdd FILL
XFILL_11_NOR2X1_61 gnd vdd FILL
XFILL_21_DFFSR_270 gnd vdd FILL
XFILL_52_DFFSR_94 gnd vdd FILL
XFILL_11_NOR2X1_72 gnd vdd FILL
XFILL_11_NOR2X1_83 gnd vdd FILL
XFILL_2_INVX1_210 gnd vdd FILL
XFILL_11_NOR2X1_94 gnd vdd FILL
XFILL_1_DFFSR_1 gnd vdd FILL
XFILL_2_INVX1_221 gnd vdd FILL
XFILL_21_DFFSR_60 gnd vdd FILL
XFILL_22_MUX2X1_14 gnd vdd FILL
XFILL_22_MUX2X1_25 gnd vdd FILL
XFILL_21_DFFSR_71 gnd vdd FILL
XFILL_6_INVX1_220 gnd vdd FILL
XFILL_22_MUX2X1_36 gnd vdd FILL
XFILL_21_DFFSR_82 gnd vdd FILL
XFILL_58_4_0 gnd vdd FILL
XFILL_21_DFFSR_93 gnd vdd FILL
XFILL_22_MUX2X1_47 gnd vdd FILL
XFILL_22_MUX2X1_58 gnd vdd FILL
XFILL_6_NOR3X1_4 gnd vdd FILL
XFILL_22_MUX2X1_69 gnd vdd FILL
XFILL_5_OAI22X1_19 gnd vdd FILL
XFILL_5_1_2 gnd vdd FILL
XFILL_52_DFFSR_180 gnd vdd FILL
XFILL_52_DFFSR_191 gnd vdd FILL
XFILL_61_DFFSR_70 gnd vdd FILL
XFILL_61_DFFSR_81 gnd vdd FILL
XFILL_61_DFFSR_92 gnd vdd FILL
XFILL_4_NAND3X1_40 gnd vdd FILL
XFILL_4_NAND3X1_51 gnd vdd FILL
XFILL_4_NAND3X1_62 gnd vdd FILL
XFILL_4_NAND3X1_73 gnd vdd FILL
XFILL_8_NAND2X1_20 gnd vdd FILL
XFILL_36_DFFSR_3 gnd vdd FILL
XFILL_4_NAND3X1_84 gnd vdd FILL
XFILL_56_DFFSR_190 gnd vdd FILL
XFILL_8_NAND2X1_31 gnd vdd FILL
XFILL_30_DFFSR_104 gnd vdd FILL
XFILL_8_NAND2X1_42 gnd vdd FILL
XFILL_4_DFFSR_50 gnd vdd FILL
XFILL_4_NAND3X1_95 gnd vdd FILL
XFILL_8_NAND2X1_53 gnd vdd FILL
XFILL_30_DFFSR_115 gnd vdd FILL
XFILL_4_DFFSR_61 gnd vdd FILL
XFILL_30_DFFSR_126 gnd vdd FILL
XFILL_8_NAND2X1_64 gnd vdd FILL
XFILL_4_DFFSR_72 gnd vdd FILL
XFILL_4_DFFSR_83 gnd vdd FILL
XFILL_30_DFFSR_137 gnd vdd FILL
XFILL_41_3_0 gnd vdd FILL
XFILL_8_NAND2X1_75 gnd vdd FILL
XFILL_30_DFFSR_148 gnd vdd FILL
XFILL_4_DFFSR_94 gnd vdd FILL
XFILL_13_0_2 gnd vdd FILL
XFILL_8_NAND2X1_86 gnd vdd FILL
XFILL_30_DFFSR_80 gnd vdd FILL
XFILL_30_DFFSR_159 gnd vdd FILL
XFILL_30_DFFSR_91 gnd vdd FILL
XFILL_34_DFFSR_103 gnd vdd FILL
XFILL_34_DFFSR_114 gnd vdd FILL
XFILL_11_NAND2X1_5 gnd vdd FILL
XFILL_16_CLKBUF1_17 gnd vdd FILL
XFILL_16_CLKBUF1_28 gnd vdd FILL
XFILL_34_DFFSR_125 gnd vdd FILL
XFILL_34_DFFSR_136 gnd vdd FILL
XFILL_16_CLKBUF1_39 gnd vdd FILL
XFILL_3_DFFSR_160 gnd vdd FILL
XFILL_11_AOI21X1_14 gnd vdd FILL
XFILL_34_DFFSR_147 gnd vdd FILL
XFILL_34_DFFSR_158 gnd vdd FILL
XFILL_11_AOI21X1_25 gnd vdd FILL
XFILL_3_DFFSR_171 gnd vdd FILL
XFILL_70_DFFSR_90 gnd vdd FILL
XFILL_11_AOI21X1_36 gnd vdd FILL
XFILL_34_DFFSR_169 gnd vdd FILL
XFILL_3_DFFSR_182 gnd vdd FILL
XFILL_3_DFFSR_193 gnd vdd FILL
XAND2X2_5 AND2X2_6/A AND2X2_5/B gnd AND2X2_5/Y vdd AND2X2
XFILL_11_AOI21X1_47 gnd vdd FILL
XFILL_38_DFFSR_102 gnd vdd FILL
XFILL_11_AOI21X1_58 gnd vdd FILL
XFILL_20_DFFSR_9 gnd vdd FILL
XFILL_11_AOI21X1_69 gnd vdd FILL
XFILL_38_DFFSR_113 gnd vdd FILL
XFILL_38_DFFSR_124 gnd vdd FILL
XFILL_38_DFFSR_135 gnd vdd FILL
XFILL_38_DFFSR_146 gnd vdd FILL
XFILL_38_DFFSR_157 gnd vdd FILL
XFILL_7_DFFSR_170 gnd vdd FILL
XFILL_58_DFFSR_7 gnd vdd FILL
XFILL_38_DFFSR_168 gnd vdd FILL
XFILL_7_DFFSR_181 gnd vdd FILL
XFILL_38_DFFSR_179 gnd vdd FILL
XFILL_11_MUX2X1_90 gnd vdd FILL
XFILL_7_DFFSR_192 gnd vdd FILL
XFILL_30_NOR3X1_15 gnd vdd FILL
XFILL_30_NOR3X1_26 gnd vdd FILL
XFILL_30_NOR3X1_37 gnd vdd FILL
XFILL_30_NOR3X1_48 gnd vdd FILL
XFILL_80_DFFSR_204 gnd vdd FILL
XFILL_80_DFFSR_215 gnd vdd FILL
XFILL_80_DFFSR_226 gnd vdd FILL
XFILL_2_5 gnd vdd FILL
XFILL_80_DFFSR_237 gnd vdd FILL
XFILL_80_DFFSR_248 gnd vdd FILL
XFILL_80_DFFSR_259 gnd vdd FILL
XFILL_49_4_0 gnd vdd FILL
XFILL_84_DFFSR_203 gnd vdd FILL
XFILL_23_CLKBUF1_30 gnd vdd FILL
XFILL_23_CLKBUF1_41 gnd vdd FILL
XFILL_84_DFFSR_214 gnd vdd FILL
XFILL_84_DFFSR_225 gnd vdd FILL
XFILL_84_DFFSR_236 gnd vdd FILL
XFILL_84_DFFSR_247 gnd vdd FILL
XFILL_6_CLKBUF1_12 gnd vdd FILL
XFILL_84_DFFSR_258 gnd vdd FILL
XFILL_84_DFFSR_269 gnd vdd FILL
XFILL_6_CLKBUF1_23 gnd vdd FILL
XFILL_44_5 gnd vdd FILL
XFILL_6_CLKBUF1_34 gnd vdd FILL
XFILL_0_INVX1_120 gnd vdd FILL
XFILL_0_INVX1_131 gnd vdd FILL
XFILL_14_MUX2X1_108 gnd vdd FILL
XFILL_14_MUX2X1_119 gnd vdd FILL
XFILL_1_AOI21X1_20 gnd vdd FILL
XFILL_0_INVX1_142 gnd vdd FILL
XFILL_0_INVX1_153 gnd vdd FILL
XFILL_1_AOI21X1_31 gnd vdd FILL
XFILL_0_INVX1_164 gnd vdd FILL
XFILL_15_AOI21X1_9 gnd vdd FILL
XFILL_1_AOI21X1_42 gnd vdd FILL
XFILL_0_INVX1_175 gnd vdd FILL
XFILL_1_AOI21X1_53 gnd vdd FILL
XFILL_0_INVX1_186 gnd vdd FILL
XFILL_11_OAI22X1_11 gnd vdd FILL
XFILL_11_OAI22X1_22 gnd vdd FILL
XFILL_1_AOI21X1_64 gnd vdd FILL
XFILL_0_INVX1_197 gnd vdd FILL
XFILL_23_DFFSR_190 gnd vdd FILL
XFILL_1_AOI21X1_75 gnd vdd FILL
XFILL_11_OAI22X1_33 gnd vdd FILL
XFILL_32_3_0 gnd vdd FILL
XFILL_11_OAI22X1_44 gnd vdd FILL
XFILL_4_INVX1_130 gnd vdd FILL
XFILL_15_OAI21X1_13 gnd vdd FILL
XFILL_4_INVX1_141 gnd vdd FILL
XFILL_4_INVX1_152 gnd vdd FILL
XFILL_15_OAI21X1_24 gnd vdd FILL
XFILL_4_NOR2X1_130 gnd vdd FILL
XFILL_4_NOR2X1_141 gnd vdd FILL
XFILL_15_OAI21X1_35 gnd vdd FILL
XFILL_4_INVX1_163 gnd vdd FILL
XFILL_15_OAI21X1_46 gnd vdd FILL
XFILL_4_INVX1_174 gnd vdd FILL
XFILL_4_INVX1_185 gnd vdd FILL
XFILL_4_NOR2X1_152 gnd vdd FILL
XFILL_4_NOR2X1_163 gnd vdd FILL
XFILL_4_NOR2X1_174 gnd vdd FILL
XFILL_4_INVX1_196 gnd vdd FILL
XFILL_4_NOR2X1_185 gnd vdd FILL
XFILL_4_NOR2X1_196 gnd vdd FILL
XFILL_21_MUX2X1_110 gnd vdd FILL
XFILL_21_MUX2X1_121 gnd vdd FILL
XFILL_2_OAI22X1_3 gnd vdd FILL
XFILL_21_MUX2X1_132 gnd vdd FILL
XFILL_21_MUX2X1_143 gnd vdd FILL
XFILL_21_MUX2X1_154 gnd vdd FILL
XFILL_21_MUX2X1_165 gnd vdd FILL
XFILL_60_13 gnd vdd FILL
XFILL_4_MUX2X1_103 gnd vdd FILL
XFILL_21_MUX2X1_176 gnd vdd FILL
XFILL_4_MUX2X1_114 gnd vdd FILL
XFILL_21_MUX2X1_187 gnd vdd FILL
XFILL_4_MUX2X1_125 gnd vdd FILL
XFILL_4_MUX2X1_136 gnd vdd FILL
XFILL_6_OAI22X1_2 gnd vdd FILL
XFILL_4_MUX2X1_147 gnd vdd FILL
XFILL_4_MUX2X1_158 gnd vdd FILL
XFILL_4_MUX2X1_169 gnd vdd FILL
XFILL_1_OAI22X1_50 gnd vdd FILL
XFILL_5_OAI21X1_30 gnd vdd FILL
XFILL_51_DFFSR_203 gnd vdd FILL
XFILL_5_OAI21X1_41 gnd vdd FILL
XFILL_51_DFFSR_214 gnd vdd FILL
XFILL_51_DFFSR_225 gnd vdd FILL
XFILL_51_DFFSR_236 gnd vdd FILL
XFILL_51_DFFSR_247 gnd vdd FILL
XFILL_51_DFFSR_258 gnd vdd FILL
XFILL_51_DFFSR_269 gnd vdd FILL
XFILL_5_DFFSR_2 gnd vdd FILL
XFILL_55_DFFSR_202 gnd vdd FILL
XFILL_55_DFFSR_213 gnd vdd FILL
XFILL_55_DFFSR_224 gnd vdd FILL
XFILL_23_3_0 gnd vdd FILL
XFILL_55_DFFSR_235 gnd vdd FILL
XFILL_75_DFFSR_1 gnd vdd FILL
XFILL_11_NAND3X1_104 gnd vdd FILL
XFILL_9_BUFX4_10 gnd vdd FILL
XFILL_55_DFFSR_246 gnd vdd FILL
XFILL_11_NAND3X1_115 gnd vdd FILL
XFILL_9_BUFX4_21 gnd vdd FILL
XFILL_55_DFFSR_257 gnd vdd FILL
XFILL_9_BUFX4_32 gnd vdd FILL
XFILL_11_NAND3X1_126 gnd vdd FILL
XFILL_55_DFFSR_268 gnd vdd FILL
XFILL_9_BUFX4_43 gnd vdd FILL
XFILL_10_CLKBUF1_9 gnd vdd FILL
XFILL_59_DFFSR_201 gnd vdd FILL
XFILL_82_DFFSR_102 gnd vdd FILL
XFILL_9_BUFX4_54 gnd vdd FILL
XFILL_44_DFFSR_19 gnd vdd FILL
XFILL_9_BUFX4_65 gnd vdd FILL
XFILL_59_DFFSR_212 gnd vdd FILL
XFILL_82_DFFSR_113 gnd vdd FILL
XFILL_82_DFFSR_124 gnd vdd FILL
XFILL_0_BUFX2_8 gnd vdd FILL
XFILL_9_BUFX4_76 gnd vdd FILL
XFILL_82_DFFSR_135 gnd vdd FILL
XFILL_59_DFFSR_223 gnd vdd FILL
XFILL_9_BUFX4_87 gnd vdd FILL
XFILL_59_DFFSR_234 gnd vdd FILL
XFILL_9_BUFX4_98 gnd vdd FILL
XFILL_82_DFFSR_146 gnd vdd FILL
XFILL_59_DFFSR_245 gnd vdd FILL
XFILL_82_DFFSR_157 gnd vdd FILL
XFILL_59_DFFSR_256 gnd vdd FILL
XFILL_59_DFFSR_267 gnd vdd FILL
XFILL_82_DFFSR_168 gnd vdd FILL
XFILL_82_DFFSR_179 gnd vdd FILL
XFILL_14_CLKBUF1_8 gnd vdd FILL
XFILL_2_DFFSR_205 gnd vdd FILL
XFILL_86_DFFSR_101 gnd vdd FILL
XFILL_2_DFFSR_216 gnd vdd FILL
XFILL_84_DFFSR_18 gnd vdd FILL
XFILL_86_DFFSR_112 gnd vdd FILL
XFILL_7_NAND3X1_17 gnd vdd FILL
XFILL_2_DFFSR_227 gnd vdd FILL
XFILL_84_DFFSR_29 gnd vdd FILL
XFILL_86_DFFSR_123 gnd vdd FILL
XFILL_86_DFFSR_134 gnd vdd FILL
XFILL_2_DFFSR_238 gnd vdd FILL
XFILL_7_NAND3X1_28 gnd vdd FILL
XFILL_86_DFFSR_145 gnd vdd FILL
XFILL_2_DFFSR_249 gnd vdd FILL
XFILL_7_NAND3X1_39 gnd vdd FILL
XFILL_2_NAND3X1_109 gnd vdd FILL
XFILL_86_DFFSR_156 gnd vdd FILL
XFILL_13_DFFSR_18 gnd vdd FILL
XFILL_10_BUFX4_103 gnd vdd FILL
XFILL_86_DFFSR_167 gnd vdd FILL
XFILL_13_DFFSR_29 gnd vdd FILL
XFILL_18_CLKBUF1_7 gnd vdd FILL
XFILL_86_DFFSR_178 gnd vdd FILL
XFILL_86_DFFSR_189 gnd vdd FILL
XFILL_6_DFFSR_204 gnd vdd FILL
XFILL_3_NAND3X1_4 gnd vdd FILL
XFILL_6_DFFSR_215 gnd vdd FILL
XFILL_6_DFFSR_226 gnd vdd FILL
XFILL_6_DFFSR_237 gnd vdd FILL
XFILL_6_DFFSR_248 gnd vdd FILL
XFILL_6_DFFSR_259 gnd vdd FILL
XFILL_14_BUFX4_102 gnd vdd FILL
XFILL_53_DFFSR_17 gnd vdd FILL
XFILL_53_DFFSR_28 gnd vdd FILL
XFILL_53_DFFSR_39 gnd vdd FILL
XFILL_7_NAND3X1_3 gnd vdd FILL
XFILL_6_4_0 gnd vdd FILL
XMUX2X1_17 BUFX4_85/Y INVX1_30/Y MUX2X1_20/S gnd DFFSR_10/D vdd MUX2X1
XFILL_0_NAND2X1_19 gnd vdd FILL
XMUX2X1_28 BUFX4_63/Y INVX1_41/Y NOR2X1_16/B gnd MUX2X1_28/Y vdd MUX2X1
XMUX2X1_39 INVX1_52/Y BUFX4_77/Y NAND2X1_5/Y gnd MUX2X1_39/Y vdd MUX2X1
XFILL_22_DFFSR_16 gnd vdd FILL
XFILL_22_DFFSR_27 gnd vdd FILL
XFILL_22_DFFSR_38 gnd vdd FILL
XFILL_13_BUFX4_70 gnd vdd FILL
XFILL_22_DFFSR_49 gnd vdd FILL
XFILL_13_BUFX4_81 gnd vdd FILL
XFILL_13_BUFX4_92 gnd vdd FILL
XFILL_10_MUX2X1_150 gnd vdd FILL
XFILL_10_MUX2X1_161 gnd vdd FILL
XFILL_10_MUX2X1_172 gnd vdd FILL
XFILL_14_3_0 gnd vdd FILL
XFILL_62_DFFSR_15 gnd vdd FILL
XFILL_10_MUX2X1_183 gnd vdd FILL
XFILL_22_DFFSR_202 gnd vdd FILL
XFILL_10_MUX2X1_194 gnd vdd FILL
XFILL_62_DFFSR_26 gnd vdd FILL
XFILL_22_DFFSR_213 gnd vdd FILL
XFILL_62_DFFSR_37 gnd vdd FILL
XFILL_62_DFFSR_48 gnd vdd FILL
XFILL_22_DFFSR_224 gnd vdd FILL
XFILL_22_DFFSR_235 gnd vdd FILL
XFILL_16_9 gnd vdd FILL
XFILL_3_AOI22X1_9 gnd vdd FILL
XFILL_62_DFFSR_59 gnd vdd FILL
XFILL_22_DFFSR_246 gnd vdd FILL
XFILL_22_DFFSR_257 gnd vdd FILL
XFILL_22_DFFSR_268 gnd vdd FILL
XFILL_26_DFFSR_201 gnd vdd FILL
XFILL_3_INVX1_208 gnd vdd FILL
XFILL_26_CLKBUF1_18 gnd vdd FILL
XFILL_26_DFFSR_212 gnd vdd FILL
XFILL_3_INVX1_219 gnd vdd FILL
XDFFSR_9 DFFSR_9/Q DFFSR_9/CLK DFFSR_9/R vdd DFFSR_9/D gnd vdd DFFSR
XFILL_26_CLKBUF1_29 gnd vdd FILL
XFILL_5_DFFSR_17 gnd vdd FILL
XFILL_26_DFFSR_223 gnd vdd FILL
XFILL_5_DFFSR_28 gnd vdd FILL
XFILL_7_AOI22X1_8 gnd vdd FILL
XFILL_26_DFFSR_234 gnd vdd FILL
XFILL_31_DFFSR_14 gnd vdd FILL
XFILL_5_DFFSR_39 gnd vdd FILL
XFILL_31_DFFSR_25 gnd vdd FILL
XFILL_26_DFFSR_245 gnd vdd FILL
XFILL_26_DFFSR_256 gnd vdd FILL
XFILL_31_DFFSR_36 gnd vdd FILL
XINVX1_210 DFFSR_80/Q gnd INVX1_210/Y vdd INVX1
XFILL_26_DFFSR_267 gnd vdd FILL
XFILL_31_DFFSR_47 gnd vdd FILL
XFILL_7_INVX1_207 gnd vdd FILL
XFILL_31_DFFSR_58 gnd vdd FILL
XINVX1_221 DFFSR_64/Q gnd OAI22X1_9/A vdd INVX1
XFILL_53_DFFSR_101 gnd vdd FILL
XFILL_7_INVX1_60 gnd vdd FILL
XFILL_31_DFFSR_69 gnd vdd FILL
XFILL_7_INVX1_71 gnd vdd FILL
XFILL_53_DFFSR_112 gnd vdd FILL
XFILL_7_INVX1_218 gnd vdd FILL
XFILL_53_DFFSR_123 gnd vdd FILL
XFILL_53_DFFSR_134 gnd vdd FILL
XFILL_4_AOI21X1_19 gnd vdd FILL
XFILL_7_INVX1_82 gnd vdd FILL
XFILL_7_INVX1_93 gnd vdd FILL
XFILL_71_DFFSR_13 gnd vdd FILL
XFILL_71_DFFSR_24 gnd vdd FILL
XFILL_53_DFFSR_145 gnd vdd FILL
XFILL_53_DFFSR_156 gnd vdd FILL
XFILL_71_DFFSR_35 gnd vdd FILL
XFILL_53_DFFSR_167 gnd vdd FILL
XFILL_53_DFFSR_178 gnd vdd FILL
XFILL_71_DFFSR_46 gnd vdd FILL
XFILL_14_MUX2X1_3 gnd vdd FILL
XFILL_71_DFFSR_57 gnd vdd FILL
XFILL_57_DFFSR_100 gnd vdd FILL
XFILL_53_DFFSR_189 gnd vdd FILL
XFILL_71_DFFSR_68 gnd vdd FILL
XFILL_57_DFFSR_111 gnd vdd FILL
XFILL_71_DFFSR_79 gnd vdd FILL
XFILL_7_NOR2X1_107 gnd vdd FILL
XFILL_57_DFFSR_122 gnd vdd FILL
XFILL_7_NOR2X1_118 gnd vdd FILL
XFILL_57_DFFSR_133 gnd vdd FILL
XFILL_57_DFFSR_144 gnd vdd FILL
XFILL_7_NOR2X1_129 gnd vdd FILL
XNAND2X1_10 INVX2_1/A INVX1_205/A gnd MUX2X1_71/S vdd NAND2X1
XFILL_13_NAND3X1_20 gnd vdd FILL
XFILL_57_DFFSR_155 gnd vdd FILL
XNAND2X1_21 BUFX4_58/Y NOR2X1_31/Y gnd OAI22X1_32/D vdd NAND2X1
XNAND2X1_32 BUFX4_2/Y NOR3X1_2/Y gnd OAI22X1_48/B vdd NAND2X1
XFILL_13_NAND3X1_31 gnd vdd FILL
XFILL_57_DFFSR_166 gnd vdd FILL
XFILL_57_DFFSR_177 gnd vdd FILL
XFILL_13_NAND3X1_42 gnd vdd FILL
XNAND2X1_43 NOR2X1_8/A INVX1_122/Y gnd NAND3X1_53/B vdd NAND2X1
XFILL_0_DFFSR_104 gnd vdd FILL
XFILL_40_DFFSR_12 gnd vdd FILL
XFILL_13_NAND3X1_53 gnd vdd FILL
XFILL_57_DFFSR_188 gnd vdd FILL
XNAND2X1_54 BUFX4_88/Y NOR2X1_34/Y gnd OAI21X1_4/B vdd NAND2X1
XFILL_13_NAND3X1_64 gnd vdd FILL
XFILL_0_DFFSR_115 gnd vdd FILL
XFILL_57_DFFSR_199 gnd vdd FILL
XFILL_40_DFFSR_23 gnd vdd FILL
XFILL_5_BUFX4_80 gnd vdd FILL
XNAND2X1_65 NOR2X1_76/Y NOR2X1_75/Y gnd NOR3X1_27/C vdd NAND2X1
XFILL_0_DFFSR_126 gnd vdd FILL
XFILL_40_DFFSR_34 gnd vdd FILL
XFILL_65_7_1 gnd vdd FILL
XFILL_33_CLKBUF1_20 gnd vdd FILL
XFILL_5_BUFX4_91 gnd vdd FILL
XFILL_13_NAND3X1_75 gnd vdd FILL
XFILL_11_NOR3X1_9 gnd vdd FILL
XFILL_40_DFFSR_45 gnd vdd FILL
XNAND2X1_76 NOR2X1_12/A NOR2X1_50/Y gnd NAND3X1_11/A vdd NAND2X1
XFILL_0_DFFSR_137 gnd vdd FILL
XFILL_13_NAND3X1_86 gnd vdd FILL
XNAND2X1_87 BUFX2_8/A BUFX2_9/A gnd INVX1_139/A vdd NAND2X1
XFILL_33_CLKBUF1_31 gnd vdd FILL
XFILL_40_DFFSR_56 gnd vdd FILL
XFILL_0_DFFSR_148 gnd vdd FILL
XFILL_13_NAND3X1_97 gnd vdd FILL
XFILL_33_CLKBUF1_42 gnd vdd FILL
XFILL_64_2_0 gnd vdd FILL
XFILL_40_DFFSR_67 gnd vdd FILL
XFILL_0_DFFSR_159 gnd vdd FILL
XFILL_40_DFFSR_78 gnd vdd FILL
XFILL_42_2 gnd vdd FILL
XFILL_40_DFFSR_89 gnd vdd FILL
XFILL_80_DFFSR_11 gnd vdd FILL
XFILL_4_DFFSR_103 gnd vdd FILL
XFILL_80_DFFSR_22 gnd vdd FILL
XFILL_4_DFFSR_114 gnd vdd FILL
XFILL_80_DFFSR_33 gnd vdd FILL
XFILL_4_DFFSR_125 gnd vdd FILL
XFILL_4_DFFSR_136 gnd vdd FILL
XFILL_80_DFFSR_44 gnd vdd FILL
XFILL_80_DFFSR_55 gnd vdd FILL
XFILL_23_MUX2X1_1 gnd vdd FILL
XFILL_4_DFFSR_147 gnd vdd FILL
XFILL_4_DFFSR_158 gnd vdd FILL
XFILL_80_DFFSR_66 gnd vdd FILL
XFILL_80_DFFSR_77 gnd vdd FILL
XFILL_4_DFFSR_169 gnd vdd FILL
XFILL_80_DFFSR_88 gnd vdd FILL
XFILL_80_DFFSR_99 gnd vdd FILL
XFILL_8_DFFSR_102 gnd vdd FILL
XFILL_12_MUX2X1_11 gnd vdd FILL
XFILL_8_DFFSR_113 gnd vdd FILL
XFILL_7_NOR2X1_4 gnd vdd FILL
XFILL_8_DFFSR_124 gnd vdd FILL
XFILL_12_MUX2X1_22 gnd vdd FILL
XFILL_8_DFFSR_135 gnd vdd FILL
XFILL_12_MUX2X1_33 gnd vdd FILL
XFILL_8_DFFSR_146 gnd vdd FILL
XFILL_12_MUX2X1_44 gnd vdd FILL
XFILL_8_DFFSR_157 gnd vdd FILL
XFILL_12_MUX2X1_55 gnd vdd FILL
XFILL_12_MUX2X1_66 gnd vdd FILL
XFILL_8_DFFSR_168 gnd vdd FILL
XFILL_4_OAI22X1_16 gnd vdd FILL
XFILL_12_MUX2X1_77 gnd vdd FILL
XFILL_8_DFFSR_179 gnd vdd FILL
XFILL_0_NOR3X1_15 gnd vdd FILL
XFILL_4_OAI22X1_27 gnd vdd FILL
XFILL_20_NOR3X1_7 gnd vdd FILL
XFILL_12_MUX2X1_88 gnd vdd FILL
XFILL_4_OAI22X1_38 gnd vdd FILL
XFILL_0_NOR3X1_26 gnd vdd FILL
XFILL_4_OAI22X1_49 gnd vdd FILL
XFILL_12_MUX2X1_99 gnd vdd FILL
XFILL_16_MUX2X1_10 gnd vdd FILL
XFILL_0_NOR3X1_37 gnd vdd FILL
XFILL_16_MUX2X1_21 gnd vdd FILL
XFILL_8_OAI21X1_18 gnd vdd FILL
XFILL_0_NOR3X1_48 gnd vdd FILL
XFILL_8_OAI21X1_29 gnd vdd FILL
XFILL_16_MUX2X1_32 gnd vdd FILL
XFILL_16_MUX2X1_43 gnd vdd FILL
XFILL_16_MUX2X1_54 gnd vdd FILL
XFILL_6_MUX2X1_2 gnd vdd FILL
XFILL_16_MUX2X1_65 gnd vdd FILL
XFILL_4_NOR3X1_14 gnd vdd FILL
XFILL_16_MUX2X1_76 gnd vdd FILL
XFILL_16_MUX2X1_87 gnd vdd FILL
XFILL_3_NAND3X1_70 gnd vdd FILL
XFILL_16_MUX2X1_98 gnd vdd FILL
XFILL_4_NOR3X1_25 gnd vdd FILL
XFILL_41_DFFSR_4 gnd vdd FILL
XFILL_4_NOR3X1_36 gnd vdd FILL
XFILL_3_NAND3X1_81 gnd vdd FILL
XFILL_9_DFFSR_3 gnd vdd FILL
XFILL_20_DFFSR_101 gnd vdd FILL
XFILL_3_NAND3X1_92 gnd vdd FILL
XFILL_4_NOR3X1_47 gnd vdd FILL
XFILL_7_NAND2X1_50 gnd vdd FILL
XFILL_20_DFFSR_112 gnd vdd FILL
XFILL_7_NAND2X1_61 gnd vdd FILL
XFILL_20_DFFSR_123 gnd vdd FILL
XFILL_20_DFFSR_134 gnd vdd FILL
XFILL_7_NAND2X1_72 gnd vdd FILL
XFILL_79_DFFSR_2 gnd vdd FILL
XFILL_20_DFFSR_145 gnd vdd FILL
XFILL_7_NAND2X1_83 gnd vdd FILL
XFILL_20_DFFSR_156 gnd vdd FILL
XFILL_8_NOR3X1_13 gnd vdd FILL
XFILL_7_NAND2X1_94 gnd vdd FILL
XFILL_8_NOR3X1_24 gnd vdd FILL
XFILL_20_DFFSR_167 gnd vdd FILL
XFILL_20_DFFSR_178 gnd vdd FILL
XFILL_3_NOR3X1_8 gnd vdd FILL
XFILL_1_INVX1_107 gnd vdd FILL
XFILL_8_NOR3X1_35 gnd vdd FILL
XFILL_20_DFFSR_189 gnd vdd FILL
XFILL_8_NOR3X1_46 gnd vdd FILL
XFILL_1_INVX1_118 gnd vdd FILL
XFILL_24_DFFSR_100 gnd vdd FILL
XFILL_1_INVX1_129 gnd vdd FILL
XFILL_24_DFFSR_111 gnd vdd FILL
XFILL_15_CLKBUF1_14 gnd vdd FILL
XFILL_15_CLKBUF1_25 gnd vdd FILL
XFILL_24_DFFSR_122 gnd vdd FILL
XFILL_15_CLKBUF1_36 gnd vdd FILL
XFILL_24_DFFSR_133 gnd vdd FILL
XFILL_4_BUFX2_9 gnd vdd FILL
XFILL_24_DFFSR_144 gnd vdd FILL
XFILL_10_AOI21X1_11 gnd vdd FILL
XFILL_24_DFFSR_155 gnd vdd FILL
XFILL_10_AOI21X1_22 gnd vdd FILL
XFILL_56_7_1 gnd vdd FILL
XFILL_10_AOI21X1_33 gnd vdd FILL
XFILL_24_DFFSR_166 gnd vdd FILL
XFILL_10_AOI21X1_44 gnd vdd FILL
XFILL_24_DFFSR_177 gnd vdd FILL
XFILL_5_INVX1_106 gnd vdd FILL
XFILL_24_DFFSR_188 gnd vdd FILL
XFILL_1_DFFSR_10 gnd vdd FILL
XFILL_55_2_0 gnd vdd FILL
XFILL_5_INVX1_117 gnd vdd FILL
XFILL_1_DFFSR_21 gnd vdd FILL
XFILL_10_AOI21X1_55 gnd vdd FILL
XFILL_10_AOI21X1_66 gnd vdd FILL
XFILL_5_INVX1_128 gnd vdd FILL
XFILL_28_DFFSR_110 gnd vdd FILL
XFILL_24_DFFSR_199 gnd vdd FILL
XFILL_5_INVX1_139 gnd vdd FILL
XFILL_10_AOI21X1_77 gnd vdd FILL
XFILL_28_DFFSR_121 gnd vdd FILL
XFILL_1_DFFSR_32 gnd vdd FILL
XFILL_1_DFFSR_43 gnd vdd FILL
XFILL_28_DFFSR_132 gnd vdd FILL
XFILL_28_DFFSR_143 gnd vdd FILL
XFILL_1_DFFSR_54 gnd vdd FILL
XFILL_28_DFFSR_154 gnd vdd FILL
XFILL_63_DFFSR_8 gnd vdd FILL
XFILL_1_DFFSR_65 gnd vdd FILL
XFILL_1_DFFSR_76 gnd vdd FILL
XFILL_28_DFFSR_165 gnd vdd FILL
XFILL_1_DFFSR_87 gnd vdd FILL
XFILL_20_NOR3X1_12 gnd vdd FILL
XFILL_28_DFFSR_176 gnd vdd FILL
XFILL_1_DFFSR_98 gnd vdd FILL
XFILL_28_DFFSR_187 gnd vdd FILL
XFILL_28_DFFSR_198 gnd vdd FILL
XFILL_20_NOR3X1_23 gnd vdd FILL
XFILL_20_NOR3X1_34 gnd vdd FILL
XFILL_70_DFFSR_201 gnd vdd FILL
XFILL_20_NOR3X1_45 gnd vdd FILL
XFILL_70_DFFSR_212 gnd vdd FILL
XFILL_70_DFFSR_223 gnd vdd FILL
XFILL_70_DFFSR_234 gnd vdd FILL
XFILL_12_NAND3X1_105 gnd vdd FILL
XFILL_70_DFFSR_245 gnd vdd FILL
XFILL_24_NOR3X1_11 gnd vdd FILL
XFILL_12_NAND3X1_116 gnd vdd FILL
XFILL_70_DFFSR_256 gnd vdd FILL
XFILL_12_NAND3X1_127 gnd vdd FILL
XFILL_24_NOR3X1_22 gnd vdd FILL
XFILL_70_DFFSR_267 gnd vdd FILL
XFILL_24_NOR3X1_33 gnd vdd FILL
XFILL_74_DFFSR_200 gnd vdd FILL
XFILL_24_NOR3X1_44 gnd vdd FILL
XFILL_74_DFFSR_211 gnd vdd FILL
XFILL_74_DFFSR_222 gnd vdd FILL
XFILL_74_DFFSR_233 gnd vdd FILL
XFILL_74_DFFSR_244 gnd vdd FILL
XFILL_3_BUFX4_3 gnd vdd FILL
XFILL_28_NOR3X1_10 gnd vdd FILL
XFILL_74_DFFSR_255 gnd vdd FILL
XFILL_5_CLKBUF1_20 gnd vdd FILL
XFILL_74_DFFSR_266 gnd vdd FILL
XFILL_28_NOR3X1_21 gnd vdd FILL
XFILL_28_NOR3X1_32 gnd vdd FILL
XFILL_5_CLKBUF1_31 gnd vdd FILL
XFILL_5_CLKBUF1_42 gnd vdd FILL
XFILL_28_NOR3X1_43 gnd vdd FILL
XFILL_78_DFFSR_210 gnd vdd FILL
XOAI22X1_3 INVX1_85/Y OAI22X1_8/B INVX1_81/Y OAI22X1_3/D gnd OAI22X1_3/Y vdd OAI22X1
XFILL_13_MUX2X1_105 gnd vdd FILL
XFILL_13_MUX2X1_116 gnd vdd FILL
XFILL_78_DFFSR_221 gnd vdd FILL
XFILL_13_MUX2X1_127 gnd vdd FILL
XFILL_13_MUX2X1_138 gnd vdd FILL
XFILL_78_DFFSR_232 gnd vdd FILL
XFILL_78_DFFSR_243 gnd vdd FILL
XFILL_13_MUX2X1_149 gnd vdd FILL
XFILL_0_AOI21X1_50 gnd vdd FILL
XFILL_78_DFFSR_254 gnd vdd FILL
XFILL_0_AOI21X1_61 gnd vdd FILL
XFILL_78_DFFSR_265 gnd vdd FILL
XFILL_0_AOI21X1_72 gnd vdd FILL
XFILL_10_OAI22X1_30 gnd vdd FILL
XFILL_33_CLKBUF1_6 gnd vdd FILL
XFILL_10_OAI22X1_41 gnd vdd FILL
XFILL_14_OAI21X1_10 gnd vdd FILL
XFILL_14_OAI21X1_21 gnd vdd FILL
XFILL_14_OAI21X1_32 gnd vdd FILL
XFILL_14_OAI21X1_43 gnd vdd FILL
XFILL_3_NOR2X1_160 gnd vdd FILL
XFILL_3_NOR2X1_171 gnd vdd FILL
XFILL_3_NOR2X1_182 gnd vdd FILL
XFILL_2_INVX1_7 gnd vdd FILL
XFILL_3_NOR2X1_193 gnd vdd FILL
XFILL_47_7_1 gnd vdd FILL
XFILL_46_2_0 gnd vdd FILL
XFILL_20_MUX2X1_140 gnd vdd FILL
XFILL_21_7 gnd vdd FILL
XFILL_20_MUX2X1_151 gnd vdd FILL
XFILL_3_MUX2X1_100 gnd vdd FILL
XFILL_20_MUX2X1_162 gnd vdd FILL
XFILL_3_MUX2X1_111 gnd vdd FILL
XFILL_20_MUX2X1_173 gnd vdd FILL
XFILL_20_MUX2X1_184 gnd vdd FILL
XFILL_3_MUX2X1_122 gnd vdd FILL
XFILL_14_6 gnd vdd FILL
XFILL_3_MUX2X1_133 gnd vdd FILL
XFILL_30_6_1 gnd vdd FILL
XFILL_3_MUX2X1_144 gnd vdd FILL
XFILL_14_BUFX4_15 gnd vdd FILL
XFILL_3_MUX2X1_155 gnd vdd FILL
XFILL_14_BUFX4_26 gnd vdd FILL
XFILL_3_MUX2X1_166 gnd vdd FILL
XFILL_14_BUFX4_37 gnd vdd FILL
XFILL_6_INVX8_1 gnd vdd FILL
XFILL_14_BUFX4_48 gnd vdd FILL
XFILL_3_MUX2X1_177 gnd vdd FILL
XDFFSR_205 INVX1_89/A DFFSR_57/CLK BUFX4_21/Y vdd MUX2X1_76/Y gnd vdd DFFSR
XFILL_3_MUX2X1_188 gnd vdd FILL
XFILL_14_BUFX4_59 gnd vdd FILL
XDFFSR_216 INVX1_83/A CLKBUF1_4/Y DFFSR_49/R vdd MUX2X1_70/Y gnd vdd DFFSR
XDFFSR_227 INVX1_67/A CLKBUF1_26/Y DFFSR_4/R vdd MUX2X1_54/Y gnd vdd DFFSR
XFILL_41_DFFSR_200 gnd vdd FILL
XDFFSR_238 INVX1_61/A DFFSR_52/CLK DFFSR_42/R vdd MUX2X1_48/Y gnd vdd DFFSR
XFILL_41_DFFSR_211 gnd vdd FILL
XDFFSR_249 INVX1_45/A CLKBUF1_5/Y DFFSR_49/R vdd MUX2X1_32/Y gnd vdd DFFSR
XFILL_3_OAI21X1_1 gnd vdd FILL
XFILL_41_DFFSR_222 gnd vdd FILL
XFILL_41_DFFSR_233 gnd vdd FILL
XFILL_41_DFFSR_244 gnd vdd FILL
XFILL_41_DFFSR_255 gnd vdd FILL
XFILL_0_NOR2X1_70 gnd vdd FILL
XFILL_0_NOR2X1_81 gnd vdd FILL
XFILL_41_DFFSR_266 gnd vdd FILL
XFILL_0_NOR2X1_92 gnd vdd FILL
XFILL_45_DFFSR_210 gnd vdd FILL
XFILL_23_DFFSR_1 gnd vdd FILL
XFILL_45_DFFSR_221 gnd vdd FILL
XFILL_80_DFFSR_2 gnd vdd FILL
XFILL_45_DFFSR_232 gnd vdd FILL
XFILL_45_DFFSR_243 gnd vdd FILL
XFILL_45_DFFSR_254 gnd vdd FILL
XFILL_45_DFFSR_265 gnd vdd FILL
XFILL_4_NOR2X1_80 gnd vdd FILL
XFILL_4_NOR2X1_91 gnd vdd FILL
XFILL_72_DFFSR_110 gnd vdd FILL
XFILL_49_DFFSR_220 gnd vdd FILL
XFILL_72_DFFSR_121 gnd vdd FILL
XFILL_72_DFFSR_132 gnd vdd FILL
XFILL_72_DFFSR_143 gnd vdd FILL
XFILL_49_DFFSR_231 gnd vdd FILL
XFILL_49_DFFSR_242 gnd vdd FILL
XFILL_9_AND2X2_8 gnd vdd FILL
XFILL_72_DFFSR_154 gnd vdd FILL
XFILL_49_DFFSR_253 gnd vdd FILL
XFILL_38_7_1 gnd vdd FILL
XFILL_72_DFFSR_165 gnd vdd FILL
XFILL_49_DFFSR_264 gnd vdd FILL
XFILL_49_DFFSR_275 gnd vdd FILL
XFILL_72_DFFSR_176 gnd vdd FILL
XFILL_8_NOR2X1_90 gnd vdd FILL
XFILL_72_DFFSR_187 gnd vdd FILL
XFILL_72_DFFSR_198 gnd vdd FILL
XFILL_37_2_0 gnd vdd FILL
XFILL_76_DFFSR_120 gnd vdd FILL
XFILL_6_NAND3X1_14 gnd vdd FILL
XFILL_76_DFFSR_131 gnd vdd FILL
XFILL_6_NAND3X1_25 gnd vdd FILL
XFILL_76_DFFSR_142 gnd vdd FILL
XFILL_6_NAND3X1_36 gnd vdd FILL
XFILL_76_DFFSR_153 gnd vdd FILL
XFILL_6_NAND3X1_47 gnd vdd FILL
XFILL_6_NAND3X1_58 gnd vdd FILL
XFILL_76_DFFSR_164 gnd vdd FILL
XFILL_45_DFFSR_5 gnd vdd FILL
XFILL_6_NAND3X1_69 gnd vdd FILL
XFILL_76_DFFSR_175 gnd vdd FILL
XFILL_76_DFFSR_186 gnd vdd FILL
XFILL_6_BUFX4_14 gnd vdd FILL
XFILL_76_DFFSR_197 gnd vdd FILL
XFILL_6_BUFX4_25 gnd vdd FILL
XFILL_6_BUFX4_36 gnd vdd FILL
XFILL_6_BUFX4_47 gnd vdd FILL
XFILL_6_BUFX4_58 gnd vdd FILL
XFILL_6_BUFX4_69 gnd vdd FILL
XFILL_21_6_1 gnd vdd FILL
XFILL_0_NAND2X1_3 gnd vdd FILL
XFILL_20_1_0 gnd vdd FILL
XFILL_4_NAND2X1_2 gnd vdd FILL
XFILL_58_DFFSR_109 gnd vdd FILL
XFILL_67_DFFSR_9 gnd vdd FILL
XFILL_13_AND2X2_2 gnd vdd FILL
XFILL_8_NAND2X1_1 gnd vdd FILL
XFILL_12_DFFSR_210 gnd vdd FILL
XFILL_12_DFFSR_221 gnd vdd FILL
XFILL_12_DFFSR_232 gnd vdd FILL
XFILL_12_DFFSR_243 gnd vdd FILL
XFILL_12_DFFSR_254 gnd vdd FILL
XFILL_12_DFFSR_265 gnd vdd FILL
XFILL_25_CLKBUF1_15 gnd vdd FILL
XFILL_10_BUFX4_30 gnd vdd FILL
XFILL_16_DFFSR_220 gnd vdd FILL
XFILL_25_CLKBUF1_26 gnd vdd FILL
XFILL_29_7_1 gnd vdd FILL
XFILL_10_BUFX4_41 gnd vdd FILL
XFILL_4_7_1 gnd vdd FILL
XFILL_25_CLKBUF1_37 gnd vdd FILL
XFILL_0_AOI21X1_8 gnd vdd FILL
XFILL_10_BUFX4_52 gnd vdd FILL
XFILL_16_DFFSR_231 gnd vdd FILL
XFILL_16_DFFSR_242 gnd vdd FILL
XFILL_28_2_0 gnd vdd FILL
XFILL_7_BUFX4_4 gnd vdd FILL
XFILL_10_BUFX4_63 gnd vdd FILL
XFILL_16_DFFSR_253 gnd vdd FILL
XFILL_3_2_0 gnd vdd FILL
XFILL_10_BUFX4_74 gnd vdd FILL
XFILL_16_DFFSR_264 gnd vdd FILL
XFILL_8_CLKBUF1_19 gnd vdd FILL
XFILL_10_BUFX4_85 gnd vdd FILL
XFILL_16_DFFSR_275 gnd vdd FILL
XFILL_10_BUFX4_96 gnd vdd FILL
XFILL_3_AOI21X1_16 gnd vdd FILL
XFILL_43_DFFSR_120 gnd vdd FILL
XFILL_43_DFFSR_131 gnd vdd FILL
XFILL_4_AOI21X1_7 gnd vdd FILL
XFILL_43_DFFSR_142 gnd vdd FILL
XFILL_3_AOI21X1_27 gnd vdd FILL
XFILL_3_AOI21X1_38 gnd vdd FILL
XFILL_3_AOI21X1_49 gnd vdd FILL
XFILL_43_DFFSR_153 gnd vdd FILL
XFILL_43_DFFSR_164 gnd vdd FILL
XFILL_43_DFFSR_175 gnd vdd FILL
XFILL_13_OAI22X1_18 gnd vdd FILL
XOAI21X1_19 INVX1_32/Y NOR2X1_51/B OAI21X1_19/C gnd NOR2X1_81/A vdd OAI21X1
XFILL_43_DFFSR_186 gnd vdd FILL
XFILL_13_OAI22X1_29 gnd vdd FILL
XFILL_43_DFFSR_197 gnd vdd FILL
XFILL_17_MUX2X1_19 gnd vdd FILL
XFILL_6_NOR2X1_104 gnd vdd FILL
XFILL_47_DFFSR_130 gnd vdd FILL
XFILL_8_AOI21X1_6 gnd vdd FILL
XFILL_12_6_1 gnd vdd FILL
XFILL_6_NOR2X1_115 gnd vdd FILL
XFILL_6_NOR2X1_126 gnd vdd FILL
XFILL_47_DFFSR_141 gnd vdd FILL
XFILL_47_DFFSR_152 gnd vdd FILL
XFILL_11_1_0 gnd vdd FILL
XFILL_6_NOR2X1_137 gnd vdd FILL
XFILL_6_NOR2X1_148 gnd vdd FILL
XFILL_13_NAND3X1_106 gnd vdd FILL
XFILL_47_DFFSR_163 gnd vdd FILL
XFILL_6_NOR2X1_159 gnd vdd FILL
XFILL_47_DFFSR_174 gnd vdd FILL
XFILL_13_NAND3X1_117 gnd vdd FILL
XFILL_13_NAND3X1_128 gnd vdd FILL
XFILL_12_NAND3X1_50 gnd vdd FILL
XFILL_47_DFFSR_185 gnd vdd FILL
XFILL_6_INVX1_8 gnd vdd FILL
XFILL_4_INVX1_20 gnd vdd FILL
XFILL_12_NAND3X1_61 gnd vdd FILL
XFILL_47_DFFSR_196 gnd vdd FILL
XFILL_4_INVX1_31 gnd vdd FILL
XFILL_12_NAND3X1_72 gnd vdd FILL
XFILL_4_INVX1_42 gnd vdd FILL
XFILL_5_AND2X2_1 gnd vdd FILL
XFILL_4_INVX1_53 gnd vdd FILL
XFILL_12_NAND3X1_83 gnd vdd FILL
XFILL_12_NAND3X1_94 gnd vdd FILL
XFILL_4_INVX1_64 gnd vdd FILL
XFILL_4_INVX1_75 gnd vdd FILL
XFILL_13_AOI22X1_3 gnd vdd FILL
XFILL_4_INVX1_86 gnd vdd FILL
XFILL_4_INVX1_97 gnd vdd FILL
XFILL_25_DFFSR_109 gnd vdd FILL
XFILL_11_MUX2X1_7 gnd vdd FILL
XFILL_23_MUX2X1_106 gnd vdd FILL
XFILL_23_MUX2X1_117 gnd vdd FILL
XFILL_17_AOI22X1_2 gnd vdd FILL
XFILL_23_MUX2X1_128 gnd vdd FILL
XFILL_23_MUX2X1_139 gnd vdd FILL
XFILL_2_BUFX4_40 gnd vdd FILL
XFILL_2_BUFX4_51 gnd vdd FILL
XFILL_29_DFFSR_108 gnd vdd FILL
XFILL_19_DFFSR_11 gnd vdd FILL
XFILL_19_DFFSR_22 gnd vdd FILL
XFILL_29_DFFSR_119 gnd vdd FILL
XFILL_2_BUFX4_62 gnd vdd FILL
XFILL_19_DFFSR_33 gnd vdd FILL
XFILL_2_BUFX4_73 gnd vdd FILL
XFILL_19_DFFSR_44 gnd vdd FILL
XFILL_2_BUFX4_84 gnd vdd FILL
XFILL_19_DFFSR_55 gnd vdd FILL
XFILL_3_OAI22X1_13 gnd vdd FILL
XFILL_2_BUFX4_95 gnd vdd FILL
XFILL_19_DFFSR_66 gnd vdd FILL
XFILL_3_OAI22X1_24 gnd vdd FILL
XFILL_19_DFFSR_77 gnd vdd FILL
XFILL_3_OAI22X1_35 gnd vdd FILL
XFILL_3_OAI22X1_46 gnd vdd FILL
XFILL_19_DFFSR_88 gnd vdd FILL
XFILL_19_DFFSR_99 gnd vdd FILL
XFILL_59_DFFSR_10 gnd vdd FILL
XFILL_7_OAI21X1_15 gnd vdd FILL
XFILL_19_2_0 gnd vdd FILL
XFILL_59_DFFSR_21 gnd vdd FILL
XFILL_7_OAI21X1_26 gnd vdd FILL
XFILL_7_OAI21X1_37 gnd vdd FILL
XFILL_59_DFFSR_32 gnd vdd FILL
XFILL_59_DFFSR_43 gnd vdd FILL
XFILL_7_OAI21X1_48 gnd vdd FILL
XFILL_59_DFFSR_54 gnd vdd FILL
XFILL_59_DFFSR_65 gnd vdd FILL
XFILL_20_MUX2X1_5 gnd vdd FILL
XFILL_59_DFFSR_76 gnd vdd FILL
XFILL_62_5_1 gnd vdd FILL
XFILL_59_DFFSR_87 gnd vdd FILL
XFILL_59_DFFSR_98 gnd vdd FILL
XFILL_61_0_0 gnd vdd FILL
XFILL_27_DFFSR_2 gnd vdd FILL
XFILL_0_NOR2X1_204 gnd vdd FILL
XFILL_10_DFFSR_120 gnd vdd FILL
XFILL_75_DFFSR_209 gnd vdd FILL
XFILL_84_DFFSR_3 gnd vdd FILL
XFILL_10_DFFSR_131 gnd vdd FILL
XFILL_4_NOR2X1_8 gnd vdd FILL
XFILL_10_DFFSR_142 gnd vdd FILL
XFILL_6_NAND2X1_80 gnd vdd FILL
XFILL_28_DFFSR_20 gnd vdd FILL
XFILL_10_DFFSR_153 gnd vdd FILL
XFILL_6_NAND2X1_91 gnd vdd FILL
XFILL_28_DFFSR_31 gnd vdd FILL
XFILL_10_DFFSR_164 gnd vdd FILL
XFILL_10_DFFSR_175 gnd vdd FILL
XFILL_28_DFFSR_42 gnd vdd FILL
XFILL_29_NOR3X1_19 gnd vdd FILL
XFILL_10_DFFSR_186 gnd vdd FILL
XFILL_12_3 gnd vdd FILL
XFILL_28_DFFSR_53 gnd vdd FILL
XFILL_28_DFFSR_64 gnd vdd FILL
XFILL_14_CLKBUF1_11 gnd vdd FILL
XFILL_10_DFFSR_197 gnd vdd FILL
XFILL_28_DFFSR_75 gnd vdd FILL
XFILL_14_CLKBUF1_22 gnd vdd FILL
XFILL_79_DFFSR_208 gnd vdd FILL
XFILL_14_DFFSR_130 gnd vdd FILL
XFILL_79_DFFSR_219 gnd vdd FILL
XFILL_28_DFFSR_86 gnd vdd FILL
XFILL_14_CLKBUF1_33 gnd vdd FILL
XFILL_14_DFFSR_141 gnd vdd FILL
XFILL_28_DFFSR_97 gnd vdd FILL
XFILL_14_DFFSR_152 gnd vdd FILL
XFILL_68_DFFSR_30 gnd vdd FILL
XFILL_14_DFFSR_163 gnd vdd FILL
XFILL_14_DFFSR_174 gnd vdd FILL
XFILL_68_DFFSR_41 gnd vdd FILL
XFILL_3_MUX2X1_6 gnd vdd FILL
XFILL_3_CLKBUF1_6 gnd vdd FILL
XFILL_68_DFFSR_52 gnd vdd FILL
XFILL_14_DFFSR_185 gnd vdd FILL
XFILL_68_DFFSR_63 gnd vdd FILL
XFILL_14_DFFSR_196 gnd vdd FILL
XFILL_68_DFFSR_74 gnd vdd FILL
XFILL_68_DFFSR_85 gnd vdd FILL
XFILL_11_DFFSR_8 gnd vdd FILL
XFILL_18_DFFSR_140 gnd vdd FILL
XFILL_68_DFFSR_96 gnd vdd FILL
XFILL_18_DFFSR_151 gnd vdd FILL
XFILL_18_DFFSR_162 gnd vdd FILL
XFILL_49_DFFSR_6 gnd vdd FILL
XFILL_18_DFFSR_173 gnd vdd FILL
XFILL_7_CLKBUF1_5 gnd vdd FILL
XFILL_18_DFFSR_184 gnd vdd FILL
XFILL_10_NOR3X1_20 gnd vdd FILL
XFILL_18_DFFSR_195 gnd vdd FILL
XFILL_10_NOR3X1_31 gnd vdd FILL
XFILL_37_DFFSR_40 gnd vdd FILL
XFILL_10_NOR3X1_42 gnd vdd FILL
XFILL_37_DFFSR_51 gnd vdd FILL
XFILL_37_DFFSR_62 gnd vdd FILL
XFILL_60_DFFSR_220 gnd vdd FILL
XFILL_3_BUFX4_100 gnd vdd FILL
XFILL_37_DFFSR_73 gnd vdd FILL
XFILL_60_DFFSR_231 gnd vdd FILL
XFILL_37_DFFSR_84 gnd vdd FILL
XFILL_60_DFFSR_242 gnd vdd FILL
XFILL_37_DFFSR_95 gnd vdd FILL
XFILL_60_DFFSR_253 gnd vdd FILL
XFILL_60_DFFSR_264 gnd vdd FILL
XFILL_14_NOR3X1_30 gnd vdd FILL
XFILL_60_DFFSR_275 gnd vdd FILL
XFILL_14_NOR3X1_41 gnd vdd FILL
XFILL_14_NOR3X1_52 gnd vdd FILL
XFILL_77_DFFSR_50 gnd vdd FILL
XFILL_77_DFFSR_61 gnd vdd FILL
XFILL_64_DFFSR_230 gnd vdd FILL
XFILL_77_DFFSR_72 gnd vdd FILL
XFILL_77_DFFSR_83 gnd vdd FILL
XFILL_64_DFFSR_241 gnd vdd FILL
XFILL_77_DFFSR_94 gnd vdd FILL
XFILL_64_DFFSR_252 gnd vdd FILL
XFILL_64_DFFSR_263 gnd vdd FILL
XFILL_64_DFFSR_274 gnd vdd FILL
XFILL_18_NOR3X1_40 gnd vdd FILL
XFILL_12_MUX2X1_102 gnd vdd FILL
XFILL_18_NOR3X1_51 gnd vdd FILL
XFILL_53_5_1 gnd vdd FILL
XFILL_12_MUX2X1_113 gnd vdd FILL
XFILL_12_MUX2X1_124 gnd vdd FILL
XFILL_0_INVX1_90 gnd vdd FILL
XFILL_12_MUX2X1_135 gnd vdd FILL
XFILL_0_BUFX2_10 gnd vdd FILL
XFILL_12_MUX2X1_146 gnd vdd FILL
XFILL_52_0_0 gnd vdd FILL
XFILL_17_NOR3X1_2 gnd vdd FILL
XFILL_68_DFFSR_240 gnd vdd FILL
XFILL_68_DFFSR_251 gnd vdd FILL
XFILL_68_DFFSR_262 gnd vdd FILL
XFILL_46_DFFSR_60 gnd vdd FILL
XFILL_12_MUX2X1_157 gnd vdd FILL
XFILL_23_CLKBUF1_3 gnd vdd FILL
XFILL_68_DFFSR_273 gnd vdd FILL
XFILL_12_MUX2X1_168 gnd vdd FILL
XFILL_46_DFFSR_71 gnd vdd FILL
XFILL_12_MUX2X1_179 gnd vdd FILL
XFILL_46_DFFSR_82 gnd vdd FILL
XFILL_46_DFFSR_93 gnd vdd FILL
XFILL_1_NOR2X1_13 gnd vdd FILL
XFILL_42_DFFSR_209 gnd vdd FILL
XFILL_1_NOR2X1_24 gnd vdd FILL
XFILL_1_NOR2X1_35 gnd vdd FILL
XFILL_1_NOR2X1_46 gnd vdd FILL
XFILL_13_OAI21X1_40 gnd vdd FILL
XFILL_1_NOR2X1_57 gnd vdd FILL
XFILL_1_NOR2X1_68 gnd vdd FILL
XFILL_1_NOR2X1_79 gnd vdd FILL
XFILL_86_DFFSR_70 gnd vdd FILL
XFILL_27_CLKBUF1_2 gnd vdd FILL
XFILL_2_NOR2X1_190 gnd vdd FILL
XFILL_86_DFFSR_81 gnd vdd FILL
XFILL_5_NOR2X1_12 gnd vdd FILL
XFILL_86_DFFSR_92 gnd vdd FILL
XFILL_46_DFFSR_208 gnd vdd FILL
XFILL_46_DFFSR_219 gnd vdd FILL
XFILL_5_NOR2X1_23 gnd vdd FILL
XFILL_8_OAI21X1_9 gnd vdd FILL
XFILL_15_DFFSR_70 gnd vdd FILL
XFILL_5_NOR2X1_34 gnd vdd FILL
XFILL_5_NOR2X1_45 gnd vdd FILL
XFILL_5_NOR2X1_56 gnd vdd FILL
XFILL_15_DFFSR_81 gnd vdd FILL
XFILL_15_DFFSR_92 gnd vdd FILL
XFILL_5_NOR2X1_67 gnd vdd FILL
XFILL_5_NOR2X1_78 gnd vdd FILL
XFILL_5_NOR2X1_89 gnd vdd FILL
XFILL_9_NOR2X1_11 gnd vdd FILL
XFILL_73_DFFSR_108 gnd vdd FILL
XFILL_73_DFFSR_119 gnd vdd FILL
XFILL_9_NOR2X1_22 gnd vdd FILL
XFILL_9_NOR2X1_33 gnd vdd FILL
XFILL_55_DFFSR_80 gnd vdd FILL
XFILL_9_NOR2X1_44 gnd vdd FILL
XFILL_9_NOR2X1_55 gnd vdd FILL
XFILL_13_OAI22X1_6 gnd vdd FILL
XFILL_9_NOR2X1_66 gnd vdd FILL
XFILL_55_DFFSR_91 gnd vdd FILL
XFILL_9_NOR2X1_77 gnd vdd FILL
XFILL_9_NOR2X1_88 gnd vdd FILL
XFILL_77_DFFSR_107 gnd vdd FILL
XFILL_9_NOR2X1_99 gnd vdd FILL
XFILL_0_NOR2X1_1 gnd vdd FILL
XFILL_77_DFFSR_118 gnd vdd FILL
XFILL_2_MUX2X1_130 gnd vdd FILL
XFILL_2_MUX2X1_141 gnd vdd FILL
XFILL_77_DFFSR_129 gnd vdd FILL
XFILL_2_MUX2X1_152 gnd vdd FILL
XFILL_2_MUX2X1_163 gnd vdd FILL
XFILL_15_NAND3X1_16 gnd vdd FILL
XFILL_17_OAI22X1_5 gnd vdd FILL
XFILL_2_MUX2X1_174 gnd vdd FILL
XFILL_15_NAND3X1_27 gnd vdd FILL
XFILL_2_MUX2X1_185 gnd vdd FILL
XFILL_15_NAND3X1_38 gnd vdd FILL
XFILL_15_NAND3X1_49 gnd vdd FILL
XFILL_24_DFFSR_90 gnd vdd FILL
XFILL_9_NOR3X1_1 gnd vdd FILL
XFILL_35_CLKBUF1_16 gnd vdd FILL
XFILL_35_CLKBUF1_27 gnd vdd FILL
XFILL_7_BUFX2_1 gnd vdd FILL
XFILL_35_CLKBUF1_38 gnd vdd FILL
XFILL_31_DFFSR_230 gnd vdd FILL
XFILL_31_DFFSR_241 gnd vdd FILL
XFILL_31_DFFSR_252 gnd vdd FILL
XFILL_44_5_1 gnd vdd FILL
XFILL_31_DFFSR_263 gnd vdd FILL
XFILL_31_DFFSR_274 gnd vdd FILL
XFILL_43_0_0 gnd vdd FILL
XFILL_35_DFFSR_240 gnd vdd FILL
XFILL_35_DFFSR_251 gnd vdd FILL
XFILL_11_BUFX4_19 gnd vdd FILL
XFILL_35_DFFSR_262 gnd vdd FILL
XFILL_35_DFFSR_273 gnd vdd FILL
XFILL_1_MUX2X1_20 gnd vdd FILL
XFILL_7_DFFSR_80 gnd vdd FILL
XFILL_1_MUX2X1_31 gnd vdd FILL
XFILL_1_MUX2X1_42 gnd vdd FILL
XFILL_7_DFFSR_91 gnd vdd FILL
XFILL_1_MUX2X1_53 gnd vdd FILL
XFILL_62_DFFSR_140 gnd vdd FILL
XFILL_1_MUX2X1_64 gnd vdd FILL
XFILL_1_MUX2X1_75 gnd vdd FILL
XFILL_62_DFFSR_151 gnd vdd FILL
XFILL_1_MUX2X1_86 gnd vdd FILL
XFILL_14_NAND3X1_107 gnd vdd FILL
XFILL_39_DFFSR_250 gnd vdd FILL
XFILL_62_DFFSR_162 gnd vdd FILL
XFILL_1_MUX2X1_97 gnd vdd FILL
XFILL_14_NAND3X1_118 gnd vdd FILL
XFILL_39_DFFSR_261 gnd vdd FILL
XFILL_39_DFFSR_272 gnd vdd FILL
XFILL_62_DFFSR_173 gnd vdd FILL
XFILL_62_DFFSR_184 gnd vdd FILL
XFILL_14_NAND3X1_129 gnd vdd FILL
XFILL_5_MUX2X1_30 gnd vdd FILL
XFILL_62_DFFSR_195 gnd vdd FILL
XFILL_13_DFFSR_208 gnd vdd FILL
XFILL_5_MUX2X1_41 gnd vdd FILL
XFILL_5_MUX2X1_52 gnd vdd FILL
XFILL_5_NAND3X1_11 gnd vdd FILL
XFILL_10_NAND3X1_8 gnd vdd FILL
XFILL_5_NAND3X1_22 gnd vdd FILL
XFILL_13_DFFSR_219 gnd vdd FILL
XFILL_5_MUX2X1_63 gnd vdd FILL
XFILL_5_NAND3X1_33 gnd vdd FILL
XFILL_66_DFFSR_150 gnd vdd FILL
XFILL_5_NAND3X1_44 gnd vdd FILL
XFILL_5_MUX2X1_74 gnd vdd FILL
XFILL_66_DFFSR_161 gnd vdd FILL
XFILL_5_MUX2X1_85 gnd vdd FILL
XFILL_5_NAND3X1_55 gnd vdd FILL
XFILL_5_MUX2X1_96 gnd vdd FILL
XFILL_50_DFFSR_6 gnd vdd FILL
XFILL_9_NAND2X1_13 gnd vdd FILL
XFILL_5_NAND3X1_66 gnd vdd FILL
XFILL_66_DFFSR_172 gnd vdd FILL
XFILL_9_NAND2X1_24 gnd vdd FILL
XFILL_5_NAND3X1_77 gnd vdd FILL
XFILL_66_DFFSR_183 gnd vdd FILL
XFILL_5_NAND3X1_88 gnd vdd FILL
XFILL_66_DFFSR_194 gnd vdd FILL
XFILL_9_NAND2X1_35 gnd vdd FILL
XFILL_17_DFFSR_207 gnd vdd FILL
XFILL_40_DFFSR_108 gnd vdd FILL
XFILL_5_NAND3X1_99 gnd vdd FILL
XFILL_9_MUX2X1_40 gnd vdd FILL
XFILL_9_NAND2X1_46 gnd vdd FILL
XFILL_9_NAND2X1_57 gnd vdd FILL
XFILL_9_MUX2X1_51 gnd vdd FILL
XFILL_14_NAND3X1_7 gnd vdd FILL
XFILL_40_DFFSR_119 gnd vdd FILL
XFILL_17_DFFSR_218 gnd vdd FILL
XFILL_9_MUX2X1_62 gnd vdd FILL
XFILL_9_NAND2X1_68 gnd vdd FILL
XFILL_17_DFFSR_229 gnd vdd FILL
XFILL_9_MUX2X1_73 gnd vdd FILL
XFILL_9_NAND2X1_79 gnd vdd FILL
XFILL_9_MUX2X1_84 gnd vdd FILL
XFILL_9_MUX2X1_95 gnd vdd FILL
XFILL_7_INVX2_1 gnd vdd FILL
XFILL_44_DFFSR_107 gnd vdd FILL
XFILL_67_4 gnd vdd FILL
XBUFX4_30 BUFX4_51/Y gnd DFFSR_57/R vdd BUFX4
XFILL_44_DFFSR_118 gnd vdd FILL
XBUFX4_41 BUFX4_3/Y gnd DFFSR_53/R vdd BUFX4
XFILL_44_DFFSR_129 gnd vdd FILL
XBUFX4_52 BUFX4_54/A gnd DFFSR_8/R vdd BUFX4
XFILL_12_AOI21X1_18 gnd vdd FILL
XBUFX4_63 INVX8_1/Y gnd BUFX4_63/Y vdd BUFX4
XFILL_12_AOI21X1_29 gnd vdd FILL
XBUFX4_74 INVX8_2/Y gnd BUFX4_74/Y vdd BUFX4
XBUFX4_85 INVX8_4/Y gnd BUFX4_85/Y vdd BUFX4
XBUFX4_96 INVX8_3/Y gnd BUFX4_96/Y vdd BUFX4
XFILL_48_DFFSR_106 gnd vdd FILL
XFILL_15_DFFSR_9 gnd vdd FILL
XFILL_48_DFFSR_117 gnd vdd FILL
XFILL_3_BUFX4_18 gnd vdd FILL
XFILL_48_DFFSR_128 gnd vdd FILL
XFILL_35_5_1 gnd vdd FILL
XFILL_3_BUFX4_29 gnd vdd FILL
XFILL_48_DFFSR_139 gnd vdd FILL
XFILL_21_MUX2X1_50 gnd vdd FILL
XFILL_21_MUX2X1_61 gnd vdd FILL
XFILL_34_0_0 gnd vdd FILL
XFILL_21_MUX2X1_72 gnd vdd FILL
XFILL_21_MUX2X1_83 gnd vdd FILL
XFILL_21_MUX2X1_94 gnd vdd FILL
XFILL_9_AOI22X1_11 gnd vdd FILL
XFILL_24_CLKBUF1_12 gnd vdd FILL
XFILL_24_CLKBUF1_23 gnd vdd FILL
XFILL_24_CLKBUF1_34 gnd vdd FILL
XFILL_0_NAND3X1_108 gnd vdd FILL
XFILL_0_NAND3X1_119 gnd vdd FILL
XFILL_7_CLKBUF1_16 gnd vdd FILL
XFILL_7_CLKBUF1_27 gnd vdd FILL
XFILL_10_AND2X2_6 gnd vdd FILL
XFILL_7_CLKBUF1_38 gnd vdd FILL
XFILL_2_AOI21X1_13 gnd vdd FILL
XFILL_2_AOI21X1_24 gnd vdd FILL
XFILL_33_DFFSR_150 gnd vdd FILL
XFILL_2_AOI21X1_35 gnd vdd FILL
XFILL_2_AOI21X1_46 gnd vdd FILL
XFILL_33_DFFSR_161 gnd vdd FILL
XFILL_2_AOI21X1_57 gnd vdd FILL
XFILL_2_AOI21X1_68 gnd vdd FILL
XFILL_33_DFFSR_172 gnd vdd FILL
XFILL_12_OAI22X1_15 gnd vdd FILL
XFILL_33_DFFSR_183 gnd vdd FILL
XFILL_12_OAI22X1_26 gnd vdd FILL
XFILL_69_DFFSR_19 gnd vdd FILL
XFILL_33_DFFSR_194 gnd vdd FILL
XFILL_2_AOI21X1_79 gnd vdd FILL
XFILL_12_OAI22X1_37 gnd vdd FILL
XFILL_5_NOR2X1_101 gnd vdd FILL
XFILL_12_OAI22X1_48 gnd vdd FILL
XFILL_5_NOR2X1_112 gnd vdd FILL
XFILL_5_NOR2X1_123 gnd vdd FILL
XFILL_5_NOR2X1_134 gnd vdd FILL
XFILL_37_DFFSR_160 gnd vdd FILL
XFILL_5_NOR2X1_145 gnd vdd FILL
XFILL_5_NOR2X1_156 gnd vdd FILL
XFILL_37_DFFSR_171 gnd vdd FILL
XFILL_5_NOR2X1_167 gnd vdd FILL
XFILL_37_DFFSR_182 gnd vdd FILL
XFILL_5_NOR2X1_178 gnd vdd FILL
XFILL_37_DFFSR_193 gnd vdd FILL
XFILL_11_DFFSR_107 gnd vdd FILL
XFILL_5_NOR2X1_189 gnd vdd FILL
XFILL_11_DFFSR_118 gnd vdd FILL
XFILL_11_NAND3X1_80 gnd vdd FILL
XFILL_11_DFFSR_129 gnd vdd FILL
XFILL_11_NAND3X1_91 gnd vdd FILL
XFILL_38_DFFSR_18 gnd vdd FILL
XFILL_38_DFFSR_29 gnd vdd FILL
XFILL_26_5_1 gnd vdd FILL
XFILL_1_5_1 gnd vdd FILL
XFILL_15_DFFSR_106 gnd vdd FILL
XFILL_22_MUX2X1_103 gnd vdd FILL
XFILL_15_DFFSR_117 gnd vdd FILL
XFILL_25_0_0 gnd vdd FILL
XFILL_0_0_0 gnd vdd FILL
XFILL_15_DFFSR_128 gnd vdd FILL
XFILL_22_MUX2X1_114 gnd vdd FILL
XFILL_15_DFFSR_139 gnd vdd FILL
XFILL_22_MUX2X1_125 gnd vdd FILL
XFILL_10_AOI21X1_2 gnd vdd FILL
XFILL_78_DFFSR_17 gnd vdd FILL
XFILL_78_DFFSR_28 gnd vdd FILL
XFILL_22_MUX2X1_136 gnd vdd FILL
XFILL_78_DFFSR_39 gnd vdd FILL
XFILL_22_MUX2X1_147 gnd vdd FILL
XFILL_22_MUX2X1_158 gnd vdd FILL
XFILL_83_DFFSR_250 gnd vdd FILL
XFILL_83_DFFSR_261 gnd vdd FILL
XFILL_19_DFFSR_105 gnd vdd FILL
XFILL_83_DFFSR_272 gnd vdd FILL
XFILL_22_MUX2X1_169 gnd vdd FILL
XFILL_5_MUX2X1_107 gnd vdd FILL
XFILL_5_MUX2X1_118 gnd vdd FILL
XFILL_1_INVX1_13 gnd vdd FILL
XFILL_19_DFFSR_116 gnd vdd FILL
XFILL_5_MUX2X1_129 gnd vdd FILL
XFILL_19_DFFSR_127 gnd vdd FILL
XFILL_1_INVX1_24 gnd vdd FILL
XFILL_19_DFFSR_138 gnd vdd FILL
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XFILL_19_DFFSR_149 gnd vdd FILL
XFILL_1_INVX1_35 gnd vdd FILL
XFILL_2_OAI22X1_10 gnd vdd FILL
XFILL_14_AOI21X1_1 gnd vdd FILL
XFILL_1_INVX1_46 gnd vdd FILL
XFILL_2_AND2X2_5 gnd vdd FILL
XFILL_2_OAI22X1_21 gnd vdd FILL
XFILL_1_INVX1_57 gnd vdd FILL
XFILL_2_OAI22X1_32 gnd vdd FILL
XFILL_1_INVX1_68 gnd vdd FILL
XFILL_2_OAI22X1_43 gnd vdd FILL
XFILL_11_NOR3X1_18 gnd vdd FILL
XFILL_87_DFFSR_260 gnd vdd FILL
XFILL_87_DFFSR_271 gnd vdd FILL
XFILL_47_DFFSR_16 gnd vdd FILL
XFILL_1_INVX1_79 gnd vdd FILL
XFILL_47_DFFSR_27 gnd vdd FILL
XFILL_6_OAI21X1_12 gnd vdd FILL
XFILL_11_NOR3X1_29 gnd vdd FILL
XFILL_47_DFFSR_38 gnd vdd FILL
XFILL_6_OAI21X1_23 gnd vdd FILL
XFILL_61_DFFSR_207 gnd vdd FILL
XFILL_47_DFFSR_49 gnd vdd FILL
XFILL_6_OAI21X1_34 gnd vdd FILL
XFILL_6_OAI21X1_45 gnd vdd FILL
XFILL_61_DFFSR_218 gnd vdd FILL
XFILL_61_DFFSR_229 gnd vdd FILL
XFILL_15_NOR3X1_17 gnd vdd FILL
XFILL_15_NOR3X1_28 gnd vdd FILL
XFILL_87_DFFSR_15 gnd vdd FILL
XFILL_87_DFFSR_26 gnd vdd FILL
XFILL_32_DFFSR_3 gnd vdd FILL
XFILL_87_DFFSR_37 gnd vdd FILL
XFILL_15_NOR3X1_39 gnd vdd FILL
XFILL_65_DFFSR_206 gnd vdd FILL
XFILL_87_DFFSR_48 gnd vdd FILL
XFILL_65_DFFSR_217 gnd vdd FILL
XFILL_87_DFFSR_59 gnd vdd FILL
XFILL_16_DFFSR_15 gnd vdd FILL
XFILL_16_DFFSR_26 gnd vdd FILL
XFILL_65_DFFSR_228 gnd vdd FILL
XFILL_9_6_1 gnd vdd FILL
XFILL_16_DFFSR_37 gnd vdd FILL
XFILL_65_DFFSR_239 gnd vdd FILL
XFILL_16_DFFSR_48 gnd vdd FILL
XFILL_19_NOR3X1_16 gnd vdd FILL
XFILL_8_1_0 gnd vdd FILL
XFILL_16_DFFSR_59 gnd vdd FILL
XFILL_19_NOR3X1_27 gnd vdd FILL
XFILL_19_NOR3X1_38 gnd vdd FILL
XFILL_19_NOR3X1_49 gnd vdd FILL
XFILL_69_DFFSR_205 gnd vdd FILL
XFILL_13_CLKBUF1_30 gnd vdd FILL
XFILL_69_DFFSR_216 gnd vdd FILL
XFILL_56_DFFSR_14 gnd vdd FILL
XFILL_13_CLKBUF1_41 gnd vdd FILL
XFILL_69_DFFSR_227 gnd vdd FILL
XFILL_56_DFFSR_25 gnd vdd FILL
XFILL_56_DFFSR_36 gnd vdd FILL
XFILL_69_DFFSR_238 gnd vdd FILL
XFILL_69_DFFSR_249 gnd vdd FILL
XFILL_56_DFFSR_47 gnd vdd FILL
XFILL_56_DFFSR_58 gnd vdd FILL
XFILL_56_DFFSR_69 gnd vdd FILL
XFILL_17_5_1 gnd vdd FILL
XFILL_16_0_0 gnd vdd FILL
XFILL_54_DFFSR_7 gnd vdd FILL
XFILL_25_DFFSR_13 gnd vdd FILL
XFILL_25_DFFSR_24 gnd vdd FILL
XFILL_25_DFFSR_35 gnd vdd FILL
XFILL_25_DFFSR_46 gnd vdd FILL
XFILL_11_NOR2X1_170 gnd vdd FILL
XFILL_25_DFFSR_57 gnd vdd FILL
XFILL_11_NOR2X1_181 gnd vdd FILL
XFILL_25_DFFSR_68 gnd vdd FILL
XFILL_11_NOR2X1_192 gnd vdd FILL
XFILL_25_DFFSR_79 gnd vdd FILL
XFILL_65_DFFSR_12 gnd vdd FILL
XFILL_50_DFFSR_250 gnd vdd FILL
XFILL_65_DFFSR_23 gnd vdd FILL
XFILL_50_DFFSR_261 gnd vdd FILL
XFILL_50_DFFSR_272 gnd vdd FILL
XFILL_65_DFFSR_34 gnd vdd FILL
XFILL_65_DFFSR_45 gnd vdd FILL
XFILL_65_DFFSR_56 gnd vdd FILL
XFILL_65_DFFSR_67 gnd vdd FILL
XFILL_65_DFFSR_78 gnd vdd FILL
XFILL_65_DFFSR_89 gnd vdd FILL
XFILL_15_NAND3X1_108 gnd vdd FILL
XFILL_54_DFFSR_260 gnd vdd FILL
XFILL_15_NAND3X1_119 gnd vdd FILL
XFILL_54_DFFSR_271 gnd vdd FILL
XFILL_8_DFFSR_14 gnd vdd FILL
XFILL_8_DFFSR_25 gnd vdd FILL
XFILL_11_MUX2X1_110 gnd vdd FILL
XFILL_34_DFFSR_11 gnd vdd FILL
XFILL_8_DFFSR_36 gnd vdd FILL
XFILL_34_DFFSR_22 gnd vdd FILL
XFILL_8_DFFSR_47 gnd vdd FILL
XFILL_11_MUX2X1_121 gnd vdd FILL
XFILL_8_DFFSR_58 gnd vdd FILL
XFILL_34_DFFSR_33 gnd vdd FILL
XFILL_8_DFFSR_69 gnd vdd FILL
XFILL_11_MUX2X1_132 gnd vdd FILL
XFILL_34_DFFSR_44 gnd vdd FILL
XFILL_11_MUX2X1_143 gnd vdd FILL
XFILL_34_DFFSR_55 gnd vdd FILL
XFILL_11_MUX2X1_154 gnd vdd FILL
XFILL_81_DFFSR_160 gnd vdd FILL
XFILL_34_DFFSR_66 gnd vdd FILL
XFILL_11_MUX2X1_165 gnd vdd FILL
XFILL_34_DFFSR_77 gnd vdd FILL
XFILL_58_DFFSR_270 gnd vdd FILL
XFILL_81_DFFSR_171 gnd vdd FILL
XFILL_34_DFFSR_88 gnd vdd FILL
XFILL_11_MUX2X1_176 gnd vdd FILL
XFILL_81_DFFSR_182 gnd vdd FILL
XFILL_11_MUX2X1_187 gnd vdd FILL
XFILL_34_DFFSR_99 gnd vdd FILL
XFILL_81_DFFSR_193 gnd vdd FILL
XFILL_32_DFFSR_206 gnd vdd FILL
XFILL_74_DFFSR_10 gnd vdd FILL
XFILL_74_DFFSR_21 gnd vdd FILL
XFILL_32_DFFSR_217 gnd vdd FILL
XFILL_1_DFFSR_230 gnd vdd FILL
XFILL_74_DFFSR_32 gnd vdd FILL
XFILL_74_DFFSR_43 gnd vdd FILL
XFILL_1_DFFSR_241 gnd vdd FILL
XFILL_32_DFFSR_228 gnd vdd FILL
XFILL_32_DFFSR_239 gnd vdd FILL
XFILL_1_DFFSR_252 gnd vdd FILL
XFILL_74_DFFSR_54 gnd vdd FILL
XFILL_1_DFFSR_263 gnd vdd FILL
XFILL_1_DFFSR_274 gnd vdd FILL
XFILL_74_DFFSR_65 gnd vdd FILL
XFILL_74_DFFSR_76 gnd vdd FILL
XFILL_85_DFFSR_170 gnd vdd FILL
XFILL_65_1 gnd vdd FILL
XFILL_74_DFFSR_87 gnd vdd FILL
XFILL_85_DFFSR_181 gnd vdd FILL
XFILL_74_DFFSR_98 gnd vdd FILL
XFILL_85_DFFSR_192 gnd vdd FILL
XFILL_36_DFFSR_205 gnd vdd FILL
XFILL_36_DFFSR_216 gnd vdd FILL
XFILL_36_DFFSR_227 gnd vdd FILL
XFILL_5_DFFSR_240 gnd vdd FILL
XFILL_5_DFFSR_251 gnd vdd FILL
XFILL_36_DFFSR_238 gnd vdd FILL
XFILL_36_DFFSR_249 gnd vdd FILL
XFILL_5_DFFSR_262 gnd vdd FILL
XFILL_43_DFFSR_20 gnd vdd FILL
XFILL_5_DFFSR_273 gnd vdd FILL
XFILL_43_DFFSR_31 gnd vdd FILL
XFILL_2_MUX2X1_18 gnd vdd FILL
XFILL_14_NOR3X1_6 gnd vdd FILL
XFILL_43_DFFSR_42 gnd vdd FILL
XFILL_63_DFFSR_105 gnd vdd FILL
XFILL_2_MUX2X1_29 gnd vdd FILL
XFILL_43_DFFSR_53 gnd vdd FILL
XFILL_43_DFFSR_64 gnd vdd FILL
XFILL_63_DFFSR_116 gnd vdd FILL
XFILL_63_DFFSR_127 gnd vdd FILL
XFILL_43_DFFSR_75 gnd vdd FILL
XFILL_63_DFFSR_138 gnd vdd FILL
XFILL_43_DFFSR_86 gnd vdd FILL
XFILL_63_DFFSR_149 gnd vdd FILL
XFILL_9_DFFSR_250 gnd vdd FILL
XFILL_43_DFFSR_97 gnd vdd FILL
XFILL_10_NAND3X1_104 gnd vdd FILL
XFILL_10_NAND3X1_115 gnd vdd FILL
XFILL_9_DFFSR_261 gnd vdd FILL
XFILL_9_DFFSR_272 gnd vdd FILL
XFILL_83_DFFSR_30 gnd vdd FILL
XFILL_10_NAND3X1_126 gnd vdd FILL
XFILL_50_3_1 gnd vdd FILL
XFILL_83_DFFSR_41 gnd vdd FILL
XFILL_6_MUX2X1_17 gnd vdd FILL
XFILL_67_DFFSR_104 gnd vdd FILL
XFILL_83_DFFSR_52 gnd vdd FILL
XFILL_6_MUX2X1_28 gnd vdd FILL
XFILL_83_DFFSR_63 gnd vdd FILL
XFILL_6_MUX2X1_39 gnd vdd FILL
XFILL_83_DFFSR_74 gnd vdd FILL
XFILL_67_DFFSR_115 gnd vdd FILL
XFILL_67_DFFSR_126 gnd vdd FILL
XFILL_12_DFFSR_30 gnd vdd FILL
XFILL_67_DFFSR_137 gnd vdd FILL
XFILL_83_DFFSR_85 gnd vdd FILL
XFILL_12_DFFSR_41 gnd vdd FILL
XFILL_67_DFFSR_148 gnd vdd FILL
XFILL_10_OAI21X1_5 gnd vdd FILL
XFILL_83_DFFSR_96 gnd vdd FILL
XFILL_1_MUX2X1_160 gnd vdd FILL
XFILL_12_DFFSR_52 gnd vdd FILL
XFILL_14_NAND3X1_13 gnd vdd FILL
XFILL_12_DFFSR_63 gnd vdd FILL
XFILL_1_MUX2X1_171 gnd vdd FILL
XFILL_67_DFFSR_159 gnd vdd FILL
XFILL_14_NAND3X1_24 gnd vdd FILL
XFILL_12_DFFSR_74 gnd vdd FILL
XFILL_1_MUX2X1_182 gnd vdd FILL
XFILL_14_NAND3X1_35 gnd vdd FILL
XFILL_12_DFFSR_85 gnd vdd FILL
XFILL_14_NAND3X1_46 gnd vdd FILL
XFILL_1_MUX2X1_193 gnd vdd FILL
XFILL_14_NAND3X1_57 gnd vdd FILL
XFILL_12_DFFSR_96 gnd vdd FILL
XFILL_14_NAND3X1_68 gnd vdd FILL
XFILL_34_CLKBUF1_13 gnd vdd FILL
XFILL_14_NAND3X1_79 gnd vdd FILL
XFILL_34_CLKBUF1_24 gnd vdd FILL
XFILL_23_NOR3X1_4 gnd vdd FILL
XFILL_52_DFFSR_40 gnd vdd FILL
XFILL_34_CLKBUF1_35 gnd vdd FILL
XFILL_2_AOI22X1_1 gnd vdd FILL
XFILL_14_OAI21X1_4 gnd vdd FILL
XFILL_52_DFFSR_51 gnd vdd FILL
XFILL_1_NAND3X1_109 gnd vdd FILL
XFILL_52_DFFSR_62 gnd vdd FILL
XFILL_11_NOR2X1_40 gnd vdd FILL
XFILL_11_NOR2X1_51 gnd vdd FILL
XFILL_52_DFFSR_73 gnd vdd FILL
XFILL_52_DFFSR_84 gnd vdd FILL
XFILL_11_NOR2X1_62 gnd vdd FILL
XFILL_21_DFFSR_260 gnd vdd FILL
XFILL_21_DFFSR_271 gnd vdd FILL
XFILL_52_DFFSR_95 gnd vdd FILL
XFILL_2_INVX1_200 gnd vdd FILL
XFILL_11_NOR2X1_73 gnd vdd FILL
XFILL_2_INVX1_211 gnd vdd FILL
XFILL_11_NOR2X1_84 gnd vdd FILL
XFILL_11_NOR2X1_95 gnd vdd FILL
XFILL_1_DFFSR_2 gnd vdd FILL
XFILL_2_INVX1_222 gnd vdd FILL
XFILL_71_DFFSR_1 gnd vdd FILL
XFILL_25_DFFSR_270 gnd vdd FILL
XFILL_21_DFFSR_50 gnd vdd FILL
XFILL_6_INVX1_210 gnd vdd FILL
XFILL_22_MUX2X1_15 gnd vdd FILL
XFILL_21_DFFSR_61 gnd vdd FILL
XFILL_6_INVX1_221 gnd vdd FILL
XFILL_21_DFFSR_72 gnd vdd FILL
XFILL_22_MUX2X1_26 gnd vdd FILL
XFILL_21_DFFSR_83 gnd vdd FILL
XFILL_22_MUX2X1_37 gnd vdd FILL
XFILL_22_MUX2X1_48 gnd vdd FILL
XFILL_21_DFFSR_94 gnd vdd FILL
XFILL_58_4_1 gnd vdd FILL
XFILL_22_MUX2X1_59 gnd vdd FILL
XFILL_6_NOR3X1_5 gnd vdd FILL
XFILL_52_DFFSR_170 gnd vdd FILL
XFILL_52_DFFSR_181 gnd vdd FILL
XFILL_61_DFFSR_60 gnd vdd FILL
XFILL_52_DFFSR_192 gnd vdd FILL
XFILL_61_DFFSR_71 gnd vdd FILL
XFILL_61_DFFSR_82 gnd vdd FILL
XFILL_61_DFFSR_93 gnd vdd FILL
XFILL_4_NAND3X1_30 gnd vdd FILL
XFILL_4_NAND3X1_41 gnd vdd FILL
XFILL_4_NAND3X1_52 gnd vdd FILL
XFILL_8_NAND2X1_10 gnd vdd FILL
XFILL_8_NAND2X1_21 gnd vdd FILL
XFILL_4_NAND3X1_63 gnd vdd FILL
XFILL_4_DFFSR_40 gnd vdd FILL
XFILL_56_DFFSR_180 gnd vdd FILL
XFILL_4_NAND3X1_74 gnd vdd FILL
XFILL_8_NAND2X1_32 gnd vdd FILL
XFILL_36_DFFSR_4 gnd vdd FILL
XFILL_4_NAND3X1_85 gnd vdd FILL
XFILL_56_DFFSR_191 gnd vdd FILL
XFILL_4_DFFSR_51 gnd vdd FILL
XFILL_4_NAND3X1_96 gnd vdd FILL
XFILL_30_DFFSR_105 gnd vdd FILL
XFILL_8_NAND2X1_43 gnd vdd FILL
XFILL_30_DFFSR_116 gnd vdd FILL
XFILL_4_DFFSR_62 gnd vdd FILL
XFILL_8_NAND2X1_54 gnd vdd FILL
XFILL_8_NAND2X1_65 gnd vdd FILL
XFILL_4_DFFSR_73 gnd vdd FILL
XFILL_30_DFFSR_127 gnd vdd FILL
XFILL_30_DFFSR_138 gnd vdd FILL
XFILL_4_DFFSR_84 gnd vdd FILL
XFILL_41_3_1 gnd vdd FILL
XFILL_8_NAND2X1_76 gnd vdd FILL
XFILL_4_DFFSR_95 gnd vdd FILL
XFILL_30_DFFSR_149 gnd vdd FILL
XFILL_8_NAND2X1_87 gnd vdd FILL
XFILL_30_DFFSR_70 gnd vdd FILL
XFILL_30_DFFSR_81 gnd vdd FILL
XFILL_30_DFFSR_92 gnd vdd FILL
XFILL_34_DFFSR_104 gnd vdd FILL
XFILL_16_CLKBUF1_18 gnd vdd FILL
XFILL_34_DFFSR_115 gnd vdd FILL
XFILL_11_NAND2X1_6 gnd vdd FILL
XFILL_16_CLKBUF1_29 gnd vdd FILL
XFILL_34_DFFSR_126 gnd vdd FILL
XFILL_34_DFFSR_137 gnd vdd FILL
XFILL_3_DFFSR_150 gnd vdd FILL
XFILL_3_DFFSR_161 gnd vdd FILL
XFILL_34_DFFSR_148 gnd vdd FILL
XFILL_11_AOI21X1_15 gnd vdd FILL
XFILL_34_DFFSR_159 gnd vdd FILL
XFILL_70_DFFSR_80 gnd vdd FILL
XFILL_3_DFFSR_172 gnd vdd FILL
XFILL_11_AOI21X1_26 gnd vdd FILL
XFILL_3_DFFSR_183 gnd vdd FILL
XFILL_70_DFFSR_91 gnd vdd FILL
XFILL_11_AOI21X1_37 gnd vdd FILL
XFILL_3_DFFSR_194 gnd vdd FILL
XFILL_11_AOI21X1_48 gnd vdd FILL
XAND2X2_6 AND2X2_6/A AND2X2_6/B gnd AND2X2_6/Y vdd AND2X2
XFILL_11_AOI21X1_59 gnd vdd FILL
XFILL_38_DFFSR_103 gnd vdd FILL
XFILL_38_DFFSR_114 gnd vdd FILL
XFILL_38_DFFSR_125 gnd vdd FILL
XFILL_38_DFFSR_136 gnd vdd FILL
XFILL_7_DFFSR_160 gnd vdd FILL
XFILL_38_DFFSR_147 gnd vdd FILL
XFILL_38_DFFSR_158 gnd vdd FILL
XFILL_7_DFFSR_171 gnd vdd FILL
XFILL_58_DFFSR_8 gnd vdd FILL
XFILL_11_MUX2X1_80 gnd vdd FILL
XFILL_38_DFFSR_169 gnd vdd FILL
XFILL_7_DFFSR_182 gnd vdd FILL
XFILL_30_NOR3X1_16 gnd vdd FILL
XFILL_11_MUX2X1_91 gnd vdd FILL
XFILL_7_DFFSR_193 gnd vdd FILL
XFILL_30_NOR3X1_27 gnd vdd FILL
XFILL_30_NOR3X1_38 gnd vdd FILL
XFILL_30_NOR3X1_49 gnd vdd FILL
XFILL_80_DFFSR_205 gnd vdd FILL
XFILL_80_DFFSR_216 gnd vdd FILL
XFILL_80_DFFSR_227 gnd vdd FILL
XFILL_80_DFFSR_238 gnd vdd FILL
XFILL_80_DFFSR_249 gnd vdd FILL
XFILL_15_MUX2X1_90 gnd vdd FILL
XFILL_49_4_1 gnd vdd FILL
XFILL_3_NOR3X1_50 gnd vdd FILL
XFILL_23_CLKBUF1_20 gnd vdd FILL
XFILL_84_DFFSR_204 gnd vdd FILL
XFILL_84_DFFSR_215 gnd vdd FILL
XFILL_23_CLKBUF1_31 gnd vdd FILL
XFILL_23_CLKBUF1_42 gnd vdd FILL
XFILL_84_DFFSR_226 gnd vdd FILL
XFILL_84_DFFSR_237 gnd vdd FILL
XFILL_84_DFFSR_248 gnd vdd FILL
XFILL_6_CLKBUF1_13 gnd vdd FILL
XFILL_84_DFFSR_259 gnd vdd FILL
XFILL_6_CLKBUF1_24 gnd vdd FILL
XFILL_0_INVX1_110 gnd vdd FILL
XFILL_6_CLKBUF1_35 gnd vdd FILL
XFILL_0_INVX1_121 gnd vdd FILL
XFILL_14_MUX2X1_109 gnd vdd FILL
XFILL_1_AOI21X1_10 gnd vdd FILL
XFILL_0_INVX1_132 gnd vdd FILL
XFILL_1_AOI21X1_21 gnd vdd FILL
XFILL_0_INVX1_143 gnd vdd FILL
XFILL_0_INVX1_154 gnd vdd FILL
XFILL_1_AOI21X1_32 gnd vdd FILL
XFILL_1_AOI21X1_43 gnd vdd FILL
XFILL_0_INVX1_165 gnd vdd FILL
XFILL_1_AOI21X1_54 gnd vdd FILL
XFILL_11_OAI22X1_12 gnd vdd FILL
XFILL_0_INVX1_176 gnd vdd FILL
XFILL_0_INVX1_187 gnd vdd FILL
XFILL_1_AOI21X1_65 gnd vdd FILL
XFILL_23_DFFSR_180 gnd vdd FILL
XFILL_0_INVX1_198 gnd vdd FILL
XFILL_11_OAI22X1_23 gnd vdd FILL
XFILL_1_AOI21X1_76 gnd vdd FILL
XFILL_11_OAI22X1_34 gnd vdd FILL
XFILL_23_DFFSR_191 gnd vdd FILL
XFILL_32_3_1 gnd vdd FILL
XFILL_4_INVX1_120 gnd vdd FILL
XFILL_11_OAI22X1_45 gnd vdd FILL
XFILL_4_INVX1_131 gnd vdd FILL
XFILL_15_OAI21X1_14 gnd vdd FILL
XFILL_4_INVX1_142 gnd vdd FILL
XFILL_4_INVX1_153 gnd vdd FILL
XFILL_15_OAI21X1_25 gnd vdd FILL
XFILL_4_NOR2X1_120 gnd vdd FILL
XFILL_4_INVX1_164 gnd vdd FILL
XFILL_15_OAI21X1_36 gnd vdd FILL
XFILL_4_NOR2X1_131 gnd vdd FILL
XFILL_4_NOR2X1_142 gnd vdd FILL
XFILL_4_NOR2X1_153 gnd vdd FILL
XFILL_4_INVX1_175 gnd vdd FILL
XFILL_15_OAI21X1_47 gnd vdd FILL
XFILL_4_INVX1_186 gnd vdd FILL
XFILL_4_NOR2X1_164 gnd vdd FILL
XFILL_4_INVX1_197 gnd vdd FILL
XFILL_27_DFFSR_190 gnd vdd FILL
XFILL_4_NOR2X1_175 gnd vdd FILL
XFILL_4_NOR2X1_186 gnd vdd FILL
XFILL_4_NOR2X1_197 gnd vdd FILL
XFILL_21_MUX2X1_100 gnd vdd FILL
XFILL_21_MUX2X1_111 gnd vdd FILL
XFILL_21_MUX2X1_122 gnd vdd FILL
XFILL_2_OAI22X1_4 gnd vdd FILL
XFILL_21_MUX2X1_133 gnd vdd FILL
XFILL_21_MUX2X1_144 gnd vdd FILL
XFILL_21_MUX2X1_155 gnd vdd FILL
XFILL_21_MUX2X1_166 gnd vdd FILL
XFILL_60_14 gnd vdd FILL
XFILL_4_MUX2X1_104 gnd vdd FILL
XFILL_4_MUX2X1_115 gnd vdd FILL
XFILL_21_MUX2X1_177 gnd vdd FILL
XFILL_21_MUX2X1_188 gnd vdd FILL
XFILL_4_MUX2X1_126 gnd vdd FILL
XFILL_4_MUX2X1_137 gnd vdd FILL
XFILL_6_OAI22X1_3 gnd vdd FILL
XFILL_4_MUX2X1_148 gnd vdd FILL
XFILL_4_MUX2X1_159 gnd vdd FILL
XFILL_1_OAI22X1_40 gnd vdd FILL
XFILL_1_OAI22X1_51 gnd vdd FILL
XFILL_5_OAI21X1_20 gnd vdd FILL
XFILL_5_OAI21X1_31 gnd vdd FILL
XFILL_51_DFFSR_204 gnd vdd FILL
XFILL_51_DFFSR_215 gnd vdd FILL
XFILL_5_OAI21X1_42 gnd vdd FILL
XFILL_51_DFFSR_226 gnd vdd FILL
XFILL_51_DFFSR_237 gnd vdd FILL
XFILL_51_DFFSR_248 gnd vdd FILL
XFILL_51_DFFSR_259 gnd vdd FILL
XFILL_5_DFFSR_3 gnd vdd FILL
XFILL_55_DFFSR_203 gnd vdd FILL
XFILL_18_DFFSR_1 gnd vdd FILL
XFILL_55_DFFSR_214 gnd vdd FILL
XFILL_55_DFFSR_225 gnd vdd FILL
XFILL_23_3_1 gnd vdd FILL
XFILL_75_DFFSR_2 gnd vdd FILL
XFILL_9_BUFX4_11 gnd vdd FILL
XFILL_55_DFFSR_236 gnd vdd FILL
XFILL_11_NAND3X1_105 gnd vdd FILL
XFILL_11_NAND3X1_116 gnd vdd FILL
XFILL_55_DFFSR_247 gnd vdd FILL
XFILL_9_BUFX4_22 gnd vdd FILL
XFILL_55_DFFSR_258 gnd vdd FILL
XFILL_55_DFFSR_269 gnd vdd FILL
XFILL_9_BUFX4_33 gnd vdd FILL
XFILL_11_NAND3X1_127 gnd vdd FILL
XFILL_9_BUFX4_44 gnd vdd FILL
XFILL_82_DFFSR_103 gnd vdd FILL
XFILL_9_BUFX4_55 gnd vdd FILL
XFILL_59_DFFSR_202 gnd vdd FILL
XFILL_9_BUFX4_66 gnd vdd FILL
XFILL_59_DFFSR_213 gnd vdd FILL
XFILL_82_DFFSR_114 gnd vdd FILL
XFILL_0_BUFX2_9 gnd vdd FILL
XFILL_9_BUFX4_77 gnd vdd FILL
XFILL_59_DFFSR_224 gnd vdd FILL
XFILL_82_DFFSR_125 gnd vdd FILL
XFILL_82_DFFSR_136 gnd vdd FILL
XFILL_59_DFFSR_235 gnd vdd FILL
XFILL_9_BUFX4_88 gnd vdd FILL
XFILL_9_BUFX4_99 gnd vdd FILL
XFILL_82_DFFSR_147 gnd vdd FILL
XFILL_82_DFFSR_158 gnd vdd FILL
XFILL_59_DFFSR_246 gnd vdd FILL
XFILL_59_DFFSR_257 gnd vdd FILL
XFILL_59_DFFSR_268 gnd vdd FILL
XFILL_82_DFFSR_169 gnd vdd FILL
XFILL_14_CLKBUF1_9 gnd vdd FILL
XFILL_2_DFFSR_206 gnd vdd FILL
XFILL_86_DFFSR_102 gnd vdd FILL
XFILL_2_DFFSR_217 gnd vdd FILL
XFILL_86_DFFSR_113 gnd vdd FILL
XFILL_84_DFFSR_19 gnd vdd FILL
XFILL_86_DFFSR_124 gnd vdd FILL
XFILL_7_NAND3X1_18 gnd vdd FILL
XFILL_2_DFFSR_228 gnd vdd FILL
XFILL_86_DFFSR_135 gnd vdd FILL
XFILL_7_NAND3X1_29 gnd vdd FILL
XFILL_2_DFFSR_239 gnd vdd FILL
XFILL_86_DFFSR_146 gnd vdd FILL
XFILL_86_DFFSR_157 gnd vdd FILL
XFILL_10_BUFX4_104 gnd vdd FILL
XFILL_13_DFFSR_19 gnd vdd FILL
XFILL_86_DFFSR_168 gnd vdd FILL
XFILL_86_DFFSR_179 gnd vdd FILL
XFILL_18_CLKBUF1_8 gnd vdd FILL
XFILL_6_DFFSR_205 gnd vdd FILL
XFILL_6_DFFSR_216 gnd vdd FILL
XFILL_3_NAND3X1_5 gnd vdd FILL
XFILL_6_DFFSR_227 gnd vdd FILL
XFILL_6_DFFSR_238 gnd vdd FILL
XFILL_6_DFFSR_249 gnd vdd FILL
XFILL_53_DFFSR_18 gnd vdd FILL
XFILL_14_BUFX4_103 gnd vdd FILL
XFILL_53_DFFSR_29 gnd vdd FILL
XFILL_7_NAND3X1_4 gnd vdd FILL
XFILL_6_4_1 gnd vdd FILL
XMUX2X1_18 BUFX4_63/Y INVX1_31/Y MUX2X1_20/S gnd DFFSR_11/D vdd MUX2X1
XMUX2X1_29 BUFX4_71/Y INVX1_42/Y NOR2X1_16/B gnd MUX2X1_29/Y vdd MUX2X1
XFILL_12_BUFX4_1 gnd vdd FILL
XFILL_22_DFFSR_17 gnd vdd FILL
XFILL_22_DFFSR_28 gnd vdd FILL
XFILL_13_BUFX4_60 gnd vdd FILL
XFILL_13_BUFX4_71 gnd vdd FILL
XFILL_22_DFFSR_39 gnd vdd FILL
XFILL_10_MUX2X1_140 gnd vdd FILL
XFILL_13_BUFX4_82 gnd vdd FILL
XFILL_13_BUFX4_93 gnd vdd FILL
XFILL_10_MUX2X1_151 gnd vdd FILL
XFILL_10_MUX2X1_162 gnd vdd FILL
XFILL_10_MUX2X1_173 gnd vdd FILL
XFILL_14_3_1 gnd vdd FILL
XFILL_71_DFFSR_190 gnd vdd FILL
XFILL_62_DFFSR_16 gnd vdd FILL
XFILL_10_MUX2X1_184 gnd vdd FILL
XFILL_22_DFFSR_203 gnd vdd FILL
XFILL_62_DFFSR_27 gnd vdd FILL
XFILL_62_DFFSR_38 gnd vdd FILL
XFILL_22_DFFSR_214 gnd vdd FILL
XFILL_22_DFFSR_225 gnd vdd FILL
XFILL_62_DFFSR_49 gnd vdd FILL
XFILL_22_DFFSR_236 gnd vdd FILL
XFILL_22_DFFSR_247 gnd vdd FILL
XFILL_22_DFFSR_258 gnd vdd FILL
XFILL_22_DFFSR_269 gnd vdd FILL
XFILL_3_INVX1_209 gnd vdd FILL
XFILL_26_DFFSR_202 gnd vdd FILL
XFILL_26_CLKBUF1_19 gnd vdd FILL
XFILL_26_DFFSR_213 gnd vdd FILL
XAOI22X1_1 AOI22X1_1/A AOI22X1_1/B AOI22X1_1/C OAI21X1_1/Y gnd BUFX4_60/A vdd AOI22X1
XFILL_5_DFFSR_18 gnd vdd FILL
XFILL_5_DFFSR_29 gnd vdd FILL
XFILL_26_DFFSR_224 gnd vdd FILL
XFILL_7_AOI22X1_9 gnd vdd FILL
XFILL_26_DFFSR_235 gnd vdd FILL
XFILL_31_DFFSR_15 gnd vdd FILL
XFILL_31_DFFSR_26 gnd vdd FILL
XFILL_26_DFFSR_246 gnd vdd FILL
XFILL_31_DFFSR_37 gnd vdd FILL
XFILL_26_DFFSR_257 gnd vdd FILL
XFILL_26_DFFSR_268 gnd vdd FILL
XINVX1_200 DFFSR_93/Q gnd INVX1_200/Y vdd INVX1
XFILL_31_DFFSR_48 gnd vdd FILL
XINVX1_211 DFFSR_72/Q gnd INVX1_211/Y vdd INVX1
XFILL_7_INVX1_208 gnd vdd FILL
XFILL_53_DFFSR_102 gnd vdd FILL
XFILL_7_INVX1_50 gnd vdd FILL
XFILL_31_DFFSR_59 gnd vdd FILL
XINVX1_222 DFFSR_65/Q gnd INVX1_222/Y vdd INVX1
XFILL_7_INVX1_61 gnd vdd FILL
XFILL_7_INVX1_219 gnd vdd FILL
XFILL_53_DFFSR_113 gnd vdd FILL
XFILL_7_INVX1_72 gnd vdd FILL
XFILL_53_DFFSR_124 gnd vdd FILL
XFILL_7_INVX1_83 gnd vdd FILL
XFILL_7_INVX1_94 gnd vdd FILL
XFILL_53_DFFSR_135 gnd vdd FILL
XFILL_53_DFFSR_146 gnd vdd FILL
XFILL_71_DFFSR_14 gnd vdd FILL
XFILL_53_DFFSR_157 gnd vdd FILL
XFILL_71_DFFSR_25 gnd vdd FILL
XFILL_71_DFFSR_36 gnd vdd FILL
XFILL_53_DFFSR_168 gnd vdd FILL
XFILL_71_DFFSR_47 gnd vdd FILL
XFILL_53_DFFSR_179 gnd vdd FILL
XFILL_71_DFFSR_58 gnd vdd FILL
XFILL_14_MUX2X1_4 gnd vdd FILL
XFILL_57_DFFSR_101 gnd vdd FILL
XFILL_71_DFFSR_69 gnd vdd FILL
XFILL_57_DFFSR_112 gnd vdd FILL
XFILL_7_NOR2X1_108 gnd vdd FILL
XFILL_7_NOR2X1_119 gnd vdd FILL
XFILL_57_DFFSR_123 gnd vdd FILL
XFILL_57_DFFSR_134 gnd vdd FILL
XNAND2X1_11 INVX2_1/A INVX1_160/Y gnd MUX2X1_86/S vdd NAND2X1
XFILL_57_DFFSR_145 gnd vdd FILL
XFILL_13_NAND3X1_10 gnd vdd FILL
XFILL_57_DFFSR_156 gnd vdd FILL
XFILL_13_NAND3X1_21 gnd vdd FILL
XNAND2X1_22 BUFX4_5/Y NOR2X1_31/Y gnd OAI21X1_8/B vdd NAND2X1
XFILL_57_DFFSR_167 gnd vdd FILL
XFILL_13_NAND3X1_32 gnd vdd FILL
XFILL_0_MUX2X1_190 gnd vdd FILL
XNAND2X1_33 BUFX4_104/Y NOR2X1_36/Y gnd OAI22X1_49/D vdd NAND2X1
XFILL_40_DFFSR_13 gnd vdd FILL
XFILL_57_DFFSR_178 gnd vdd FILL
XFILL_2_INVX8_1 gnd vdd FILL
XFILL_0_DFFSR_105 gnd vdd FILL
XNAND2X1_44 BUFX4_6/Y NOR3X1_2/Y gnd OAI21X1_9/B vdd NAND2X1
XFILL_13_NAND3X1_43 gnd vdd FILL
XNAND2X1_55 NOR2X1_56/Y NOR2X1_55/Y gnd NOR3X1_11/C vdd NAND2X1
XFILL_5_BUFX4_70 gnd vdd FILL
XFILL_57_DFFSR_189 gnd vdd FILL
XFILL_13_NAND3X1_54 gnd vdd FILL
XFILL_13_NAND3X1_65 gnd vdd FILL
XNAND2X1_66 NOR2X1_78/Y NOR2X1_77/Y gnd NOR3X1_27/B vdd NAND2X1
XFILL_5_BUFX4_81 gnd vdd FILL
XFILL_40_DFFSR_24 gnd vdd FILL
XFILL_0_DFFSR_116 gnd vdd FILL
XFILL_33_CLKBUF1_10 gnd vdd FILL
XFILL_33_CLKBUF1_21 gnd vdd FILL
XFILL_40_DFFSR_35 gnd vdd FILL
XFILL_13_NAND3X1_76 gnd vdd FILL
XNAND2X1_77 NOR2X1_9/A INVX1_122/Y gnd NAND3X1_11/B vdd NAND2X1
XFILL_0_DFFSR_127 gnd vdd FILL
XFILL_0_DFFSR_138 gnd vdd FILL
XFILL_65_7_2 gnd vdd FILL
XFILL_5_BUFX4_92 gnd vdd FILL
XFILL_40_DFFSR_46 gnd vdd FILL
XFILL_13_NAND3X1_87 gnd vdd FILL
XFILL_33_CLKBUF1_32 gnd vdd FILL
XFILL_0_DFFSR_149 gnd vdd FILL
XFILL_40_DFFSR_57 gnd vdd FILL
XNAND2X1_88 INVX1_136/Y INVX1_140/Y gnd NOR2X1_21/B vdd NAND2X1
XFILL_64_2_1 gnd vdd FILL
XFILL_40_DFFSR_68 gnd vdd FILL
XFILL_13_NAND3X1_98 gnd vdd FILL
XFILL_42_3 gnd vdd FILL
XFILL_40_DFFSR_79 gnd vdd FILL
XFILL_4_DFFSR_104 gnd vdd FILL
XFILL_80_DFFSR_12 gnd vdd FILL
XFILL_80_DFFSR_23 gnd vdd FILL
XFILL_4_DFFSR_115 gnd vdd FILL
XFILL_4_DFFSR_126 gnd vdd FILL
XFILL_80_DFFSR_34 gnd vdd FILL
XFILL_4_DFFSR_137 gnd vdd FILL
XFILL_23_MUX2X1_2 gnd vdd FILL
XFILL_80_DFFSR_45 gnd vdd FILL
XFILL_80_DFFSR_56 gnd vdd FILL
XFILL_4_DFFSR_148 gnd vdd FILL
XFILL_80_DFFSR_67 gnd vdd FILL
XFILL_4_DFFSR_159 gnd vdd FILL
XFILL_80_DFFSR_78 gnd vdd FILL
XFILL_28_1 gnd vdd FILL
XFILL_80_DFFSR_89 gnd vdd FILL
XFILL_8_DFFSR_103 gnd vdd FILL
XFILL_8_DFFSR_114 gnd vdd FILL
XFILL_12_MUX2X1_12 gnd vdd FILL
XFILL_7_NOR2X1_5 gnd vdd FILL
XFILL_12_MUX2X1_23 gnd vdd FILL
XFILL_8_DFFSR_125 gnd vdd FILL
XFILL_8_DFFSR_136 gnd vdd FILL
XFILL_12_MUX2X1_34 gnd vdd FILL
XFILL_12_MUX2X1_45 gnd vdd FILL
XFILL_8_DFFSR_147 gnd vdd FILL
XFILL_8_DFFSR_158 gnd vdd FILL
XFILL_12_MUX2X1_56 gnd vdd FILL
XFILL_4_OAI22X1_17 gnd vdd FILL
XFILL_8_DFFSR_169 gnd vdd FILL
XFILL_12_MUX2X1_67 gnd vdd FILL
XFILL_20_NOR3X1_8 gnd vdd FILL
XFILL_4_OAI22X1_28 gnd vdd FILL
XFILL_0_NOR3X1_16 gnd vdd FILL
XFILL_12_MUX2X1_78 gnd vdd FILL
XFILL_0_NOR3X1_27 gnd vdd FILL
XFILL_12_MUX2X1_89 gnd vdd FILL
XFILL_4_OAI22X1_39 gnd vdd FILL
XFILL_16_MUX2X1_11 gnd vdd FILL
XFILL_16_MUX2X1_22 gnd vdd FILL
XFILL_0_NOR3X1_38 gnd vdd FILL
XFILL_0_NOR3X1_49 gnd vdd FILL
XFILL_17_AOI22X1_10 gnd vdd FILL
XFILL_8_OAI21X1_19 gnd vdd FILL
XFILL_16_MUX2X1_33 gnd vdd FILL
XFILL_16_MUX2X1_44 gnd vdd FILL
XFILL_16_MUX2X1_55 gnd vdd FILL
XFILL_6_MUX2X1_3 gnd vdd FILL
XFILL_16_MUX2X1_66 gnd vdd FILL
XFILL_16_MUX2X1_77 gnd vdd FILL
XFILL_3_NAND3X1_60 gnd vdd FILL
XFILL_4_NOR3X1_15 gnd vdd FILL
XFILL_16_MUX2X1_88 gnd vdd FILL
XFILL_4_NOR3X1_26 gnd vdd FILL
XFILL_41_DFFSR_5 gnd vdd FILL
XFILL_16_MUX2X1_99 gnd vdd FILL
XFILL_3_NAND3X1_71 gnd vdd FILL
XFILL_4_NOR3X1_37 gnd vdd FILL
XFILL_9_DFFSR_4 gnd vdd FILL
XFILL_20_DFFSR_102 gnd vdd FILL
XFILL_3_NAND3X1_82 gnd vdd FILL
XFILL_7_NAND2X1_40 gnd vdd FILL
XFILL_3_NAND3X1_93 gnd vdd FILL
XFILL_4_NOR3X1_48 gnd vdd FILL
XFILL_7_NAND2X1_51 gnd vdd FILL
XFILL_20_DFFSR_113 gnd vdd FILL
XFILL_20_DFFSR_124 gnd vdd FILL
XFILL_7_NAND2X1_62 gnd vdd FILL
XFILL_7_NAND2X1_73 gnd vdd FILL
XFILL_20_DFFSR_135 gnd vdd FILL
XFILL_79_DFFSR_3 gnd vdd FILL
XFILL_20_DFFSR_146 gnd vdd FILL
XFILL_7_NAND2X1_84 gnd vdd FILL
XFILL_20_DFFSR_157 gnd vdd FILL
XFILL_8_NOR3X1_14 gnd vdd FILL
XFILL_7_NAND2X1_95 gnd vdd FILL
XFILL_3_NOR3X1_9 gnd vdd FILL
XFILL_20_DFFSR_168 gnd vdd FILL
XFILL_8_NOR3X1_25 gnd vdd FILL
XFILL_20_DFFSR_179 gnd vdd FILL
XFILL_1_INVX1_108 gnd vdd FILL
XFILL_8_NOR3X1_36 gnd vdd FILL
XFILL_24_DFFSR_101 gnd vdd FILL
XFILL_8_NOR3X1_47 gnd vdd FILL
XFILL_15_CLKBUF1_15 gnd vdd FILL
XFILL_24_DFFSR_112 gnd vdd FILL
XFILL_1_INVX1_119 gnd vdd FILL
XFILL_15_CLKBUF1_26 gnd vdd FILL
XFILL_24_DFFSR_123 gnd vdd FILL
XFILL_24_DFFSR_134 gnd vdd FILL
XFILL_15_CLKBUF1_37 gnd vdd FILL
XFILL_24_DFFSR_145 gnd vdd FILL
XFILL_10_AOI21X1_12 gnd vdd FILL
XFILL_24_DFFSR_156 gnd vdd FILL
XFILL_24_DFFSR_167 gnd vdd FILL
XFILL_10_AOI21X1_23 gnd vdd FILL
XFILL_10_AOI21X1_34 gnd vdd FILL
XFILL_56_7_2 gnd vdd FILL
XFILL_10_AOI21X1_45 gnd vdd FILL
XFILL_24_DFFSR_178 gnd vdd FILL
XFILL_5_INVX1_107 gnd vdd FILL
XFILL_1_DFFSR_11 gnd vdd FILL
XFILL_28_DFFSR_100 gnd vdd FILL
XFILL_24_DFFSR_189 gnd vdd FILL
XFILL_10_AOI21X1_56 gnd vdd FILL
XFILL_10_AOI21X1_67 gnd vdd FILL
XFILL_55_2_1 gnd vdd FILL
XFILL_5_INVX1_118 gnd vdd FILL
XFILL_1_DFFSR_22 gnd vdd FILL
XFILL_28_DFFSR_111 gnd vdd FILL
XFILL_5_INVX1_129 gnd vdd FILL
XFILL_28_DFFSR_122 gnd vdd FILL
XFILL_1_DFFSR_33 gnd vdd FILL
XFILL_10_AOI21X1_78 gnd vdd FILL
XFILL_1_DFFSR_44 gnd vdd FILL
XFILL_28_DFFSR_133 gnd vdd FILL
XFILL_1_DFFSR_55 gnd vdd FILL
XFILL_28_DFFSR_144 gnd vdd FILL
XFILL_63_DFFSR_9 gnd vdd FILL
XFILL_28_DFFSR_155 gnd vdd FILL
XFILL_1_DFFSR_66 gnd vdd FILL
XFILL_1_DFFSR_77 gnd vdd FILL
XFILL_28_DFFSR_166 gnd vdd FILL
XFILL_1_DFFSR_88 gnd vdd FILL
XFILL_28_DFFSR_177 gnd vdd FILL
XFILL_20_NOR3X1_13 gnd vdd FILL
XFILL_1_DFFSR_99 gnd vdd FILL
XFILL_20_NOR3X1_24 gnd vdd FILL
XFILL_28_DFFSR_188 gnd vdd FILL
XFILL_20_NOR3X1_35 gnd vdd FILL
XFILL_28_DFFSR_199 gnd vdd FILL
XFILL_70_DFFSR_202 gnd vdd FILL
XFILL_20_NOR3X1_46 gnd vdd FILL
XFILL_70_DFFSR_213 gnd vdd FILL
XFILL_70_DFFSR_224 gnd vdd FILL
XFILL_70_DFFSR_235 gnd vdd FILL
XFILL_12_NAND3X1_106 gnd vdd FILL
XFILL_12_NAND3X1_117 gnd vdd FILL
XFILL_70_DFFSR_246 gnd vdd FILL
XFILL_12_NAND3X1_128 gnd vdd FILL
XFILL_24_NOR3X1_12 gnd vdd FILL
XFILL_70_DFFSR_257 gnd vdd FILL
XFILL_70_DFFSR_268 gnd vdd FILL
XFILL_49_DFFSR_90 gnd vdd FILL
XFILL_24_NOR3X1_23 gnd vdd FILL
XFILL_24_NOR3X1_34 gnd vdd FILL
XFILL_24_NOR3X1_45 gnd vdd FILL
XFILL_74_DFFSR_201 gnd vdd FILL
XFILL_74_DFFSR_212 gnd vdd FILL
XFILL_74_DFFSR_223 gnd vdd FILL
XFILL_74_DFFSR_234 gnd vdd FILL
XFILL_74_DFFSR_245 gnd vdd FILL
XFILL_3_BUFX4_4 gnd vdd FILL
XFILL_28_NOR3X1_11 gnd vdd FILL
XFILL_5_CLKBUF1_10 gnd vdd FILL
XFILL_74_DFFSR_256 gnd vdd FILL
XFILL_5_CLKBUF1_21 gnd vdd FILL
XFILL_74_DFFSR_267 gnd vdd FILL
XFILL_28_NOR3X1_22 gnd vdd FILL
XFILL_5_CLKBUF1_32 gnd vdd FILL
XFILL_28_NOR3X1_33 gnd vdd FILL
XFILL_28_NOR3X1_44 gnd vdd FILL
XFILL_78_DFFSR_200 gnd vdd FILL
XFILL_13_MUX2X1_106 gnd vdd FILL
XFILL_13_MUX2X1_117 gnd vdd FILL
XFILL_78_DFFSR_211 gnd vdd FILL
XOAI22X1_4 OAI22X1_4/A OAI22X1_4/B OAI22X1_4/C OAI22X1_4/D gnd OAI22X1_4/Y vdd OAI22X1
XFILL_78_DFFSR_222 gnd vdd FILL
XFILL_78_DFFSR_233 gnd vdd FILL
XFILL_13_MUX2X1_128 gnd vdd FILL
XFILL_0_AOI21X1_40 gnd vdd FILL
XFILL_13_MUX2X1_139 gnd vdd FILL
XFILL_78_DFFSR_244 gnd vdd FILL
XFILL_0_AOI21X1_51 gnd vdd FILL
XFILL_78_DFFSR_255 gnd vdd FILL
XFILL_0_AOI21X1_62 gnd vdd FILL
XFILL_0_AOI21X1_73 gnd vdd FILL
XFILL_10_OAI22X1_20 gnd vdd FILL
XFILL_78_DFFSR_266 gnd vdd FILL
XFILL_33_CLKBUF1_7 gnd vdd FILL
XFILL_10_OAI22X1_31 gnd vdd FILL
XFILL_10_OAI22X1_42 gnd vdd FILL
XFILL_14_OAI21X1_11 gnd vdd FILL
XFILL_14_OAI21X1_22 gnd vdd FILL
XFILL_14_OAI21X1_33 gnd vdd FILL
XFILL_14_OAI21X1_44 gnd vdd FILL
XFILL_3_NOR2X1_150 gnd vdd FILL
XFILL_3_NOR2X1_161 gnd vdd FILL
XFILL_3_NOR2X1_172 gnd vdd FILL
XFILL_2_INVX1_8 gnd vdd FILL
XFILL_3_NOR2X1_183 gnd vdd FILL
XFILL_3_NOR2X1_194 gnd vdd FILL
XFILL_47_7_2 gnd vdd FILL
XFILL_46_2_1 gnd vdd FILL
XFILL_20_MUX2X1_130 gnd vdd FILL
XFILL_20_MUX2X1_141 gnd vdd FILL
XFILL_21_8 gnd vdd FILL
XFILL_20_MUX2X1_152 gnd vdd FILL
XFILL_20_MUX2X1_163 gnd vdd FILL
XFILL_3_MUX2X1_101 gnd vdd FILL
XFILL_20_MUX2X1_174 gnd vdd FILL
XFILL_3_MUX2X1_112 gnd vdd FILL
XFILL_3_MUX2X1_123 gnd vdd FILL
XFILL_20_MUX2X1_185 gnd vdd FILL
XFILL_14_7 gnd vdd FILL
XFILL_3_MUX2X1_134 gnd vdd FILL
XFILL_30_6_2 gnd vdd FILL
XFILL_3_MUX2X1_145 gnd vdd FILL
XFILL_14_BUFX4_16 gnd vdd FILL
XFILL_14_BUFX4_27 gnd vdd FILL
XFILL_3_MUX2X1_156 gnd vdd FILL
XFILL_3_MUX2X1_167 gnd vdd FILL
XFILL_14_BUFX4_38 gnd vdd FILL
XFILL_3_MUX2X1_178 gnd vdd FILL
XFILL_14_BUFX4_49 gnd vdd FILL
XFILL_3_MUX2X1_189 gnd vdd FILL
XFILL_6_INVX8_2 gnd vdd FILL
XDFFSR_206 INVX1_91/A DFFSR_45/CLK BUFX4_13/Y vdd MUX2X1_77/Y gnd vdd DFFSR
XDFFSR_217 INVX1_84/A DFFSR_45/CLK DFFSR_57/R vdd MUX2X1_71/Y gnd vdd DFFSR
XDFFSR_228 INVX1_69/A DFFSR_7/CLK DFFSR_26/R vdd MUX2X1_55/Y gnd vdd DFFSR
XFILL_41_DFFSR_201 gnd vdd FILL
XDFFSR_239 INVX1_62/A DFFSR_2/CLK BUFX4_50/Y vdd MUX2X1_49/Y gnd vdd DFFSR
XFILL_41_DFFSR_212 gnd vdd FILL
XFILL_3_OAI21X1_2 gnd vdd FILL
XFILL_4_OAI21X1_50 gnd vdd FILL
XFILL_41_DFFSR_223 gnd vdd FILL
XFILL_41_DFFSR_234 gnd vdd FILL
XFILL_0_NOR2X1_60 gnd vdd FILL
XFILL_41_DFFSR_245 gnd vdd FILL
XFILL_0_NOR2X1_71 gnd vdd FILL
XFILL_41_DFFSR_256 gnd vdd FILL
XFILL_41_DFFSR_267 gnd vdd FILL
XFILL_0_NOR2X1_82 gnd vdd FILL
XFILL_0_NOR2X1_93 gnd vdd FILL
XFILL_45_DFFSR_200 gnd vdd FILL
XFILL_45_DFFSR_211 gnd vdd FILL
XFILL_23_DFFSR_2 gnd vdd FILL
XFILL_45_DFFSR_222 gnd vdd FILL
XFILL_7_OAI21X1_1 gnd vdd FILL
XFILL_80_DFFSR_3 gnd vdd FILL
XFILL_45_DFFSR_233 gnd vdd FILL
XFILL_45_DFFSR_244 gnd vdd FILL
XFILL_45_DFFSR_255 gnd vdd FILL
XFILL_4_NOR2X1_70 gnd vdd FILL
XFILL_4_NOR2X1_81 gnd vdd FILL
XFILL_45_DFFSR_266 gnd vdd FILL
XFILL_4_NOR2X1_92 gnd vdd FILL
XFILL_72_DFFSR_100 gnd vdd FILL
XFILL_72_DFFSR_111 gnd vdd FILL
XFILL_49_DFFSR_210 gnd vdd FILL
XFILL_49_DFFSR_221 gnd vdd FILL
XFILL_72_DFFSR_122 gnd vdd FILL
XFILL_72_DFFSR_133 gnd vdd FILL
XFILL_49_DFFSR_232 gnd vdd FILL
XFILL_49_DFFSR_243 gnd vdd FILL
XFILL_72_DFFSR_144 gnd vdd FILL
XFILL_72_DFFSR_155 gnd vdd FILL
XFILL_49_DFFSR_254 gnd vdd FILL
XFILL_72_DFFSR_166 gnd vdd FILL
XFILL_38_7_2 gnd vdd FILL
XFILL_8_NOR2X1_80 gnd vdd FILL
XFILL_49_DFFSR_265 gnd vdd FILL
XFILL_72_DFFSR_177 gnd vdd FILL
XFILL_37_2_1 gnd vdd FILL
XFILL_72_DFFSR_188 gnd vdd FILL
XFILL_8_NOR2X1_91 gnd vdd FILL
XFILL_76_DFFSR_110 gnd vdd FILL
XFILL_72_DFFSR_199 gnd vdd FILL
XFILL_76_DFFSR_121 gnd vdd FILL
XFILL_6_NAND3X1_15 gnd vdd FILL
XFILL_76_DFFSR_132 gnd vdd FILL
XFILL_6_NAND3X1_26 gnd vdd FILL
XFILL_76_DFFSR_143 gnd vdd FILL
XFILL_6_NAND3X1_37 gnd vdd FILL
XFILL_76_DFFSR_154 gnd vdd FILL
XFILL_6_NAND3X1_48 gnd vdd FILL
XFILL_6_NAND3X1_59 gnd vdd FILL
XFILL_76_DFFSR_165 gnd vdd FILL
XFILL_45_DFFSR_6 gnd vdd FILL
XFILL_76_DFFSR_176 gnd vdd FILL
XFILL_6_BUFX4_15 gnd vdd FILL
XFILL_76_DFFSR_187 gnd vdd FILL
XFILL_76_DFFSR_198 gnd vdd FILL
XFILL_6_BUFX4_26 gnd vdd FILL
XFILL_6_BUFX4_37 gnd vdd FILL
XFILL_6_BUFX4_48 gnd vdd FILL
XFILL_6_BUFX4_59 gnd vdd FILL
XFILL_21_6_2 gnd vdd FILL
XFILL_0_NAND2X1_4 gnd vdd FILL
XFILL_20_1_1 gnd vdd FILL
XFILL_4_NAND2X1_3 gnd vdd FILL
XFILL_13_AND2X2_3 gnd vdd FILL
XFILL_8_NAND2X1_2 gnd vdd FILL
XFILL_12_DFFSR_200 gnd vdd FILL
XFILL_12_DFFSR_211 gnd vdd FILL
XFILL_12_DFFSR_222 gnd vdd FILL
XFILL_12_DFFSR_233 gnd vdd FILL
XFILL_12_DFFSR_244 gnd vdd FILL
XFILL_12_DFFSR_255 gnd vdd FILL
XFILL_12_DFFSR_266 gnd vdd FILL
XFILL_10_BUFX4_20 gnd vdd FILL
XFILL_25_CLKBUF1_16 gnd vdd FILL
XFILL_16_DFFSR_210 gnd vdd FILL
XFILL_25_CLKBUF1_27 gnd vdd FILL
XFILL_10_BUFX4_31 gnd vdd FILL
XFILL_16_DFFSR_221 gnd vdd FILL
XFILL_29_7_2 gnd vdd FILL
XFILL_25_CLKBUF1_38 gnd vdd FILL
XFILL_0_AOI21X1_9 gnd vdd FILL
XFILL_10_BUFX4_42 gnd vdd FILL
XFILL_4_7_2 gnd vdd FILL
XFILL_16_DFFSR_232 gnd vdd FILL
XFILL_10_BUFX4_53 gnd vdd FILL
XFILL_16_DFFSR_243 gnd vdd FILL
XFILL_10_BUFX4_64 gnd vdd FILL
XFILL_3_2_1 gnd vdd FILL
XFILL_28_2_1 gnd vdd FILL
XFILL_16_DFFSR_254 gnd vdd FILL
XFILL_7_BUFX4_5 gnd vdd FILL
XFILL_16_DFFSR_265 gnd vdd FILL
XFILL_10_BUFX4_75 gnd vdd FILL
XFILL_10_BUFX4_86 gnd vdd FILL
XFILL_10_BUFX4_97 gnd vdd FILL
XFILL_43_DFFSR_110 gnd vdd FILL
XFILL_3_AOI21X1_17 gnd vdd FILL
XFILL_43_DFFSR_121 gnd vdd FILL
XFILL_43_DFFSR_132 gnd vdd FILL
XFILL_4_AOI21X1_8 gnd vdd FILL
XFILL_3_AOI21X1_28 gnd vdd FILL
XFILL_43_DFFSR_143 gnd vdd FILL
XFILL_43_DFFSR_154 gnd vdd FILL
XFILL_3_AOI21X1_39 gnd vdd FILL
XFILL_43_DFFSR_165 gnd vdd FILL
XFILL_13_OAI22X1_19 gnd vdd FILL
XFILL_43_DFFSR_176 gnd vdd FILL
XFILL_43_DFFSR_187 gnd vdd FILL
XFILL_43_DFFSR_198 gnd vdd FILL
XFILL_6_NOR2X1_105 gnd vdd FILL
XFILL_47_DFFSR_120 gnd vdd FILL
XFILL_6_NOR2X1_116 gnd vdd FILL
XFILL_12_6_2 gnd vdd FILL
XFILL_47_DFFSR_131 gnd vdd FILL
XFILL_8_AOI21X1_7 gnd vdd FILL
XFILL_47_DFFSR_142 gnd vdd FILL
XFILL_6_NOR2X1_127 gnd vdd FILL
XFILL_47_DFFSR_153 gnd vdd FILL
XFILL_11_1_1 gnd vdd FILL
XFILL_6_NOR2X1_138 gnd vdd FILL
XFILL_6_NOR2X1_149 gnd vdd FILL
XFILL_13_NAND3X1_107 gnd vdd FILL
XFILL_47_DFFSR_164 gnd vdd FILL
XFILL_47_DFFSR_175 gnd vdd FILL
XFILL_13_NAND3X1_118 gnd vdd FILL
XFILL_12_NAND3X1_40 gnd vdd FILL
XFILL_6_INVX1_9 gnd vdd FILL
XFILL_13_NAND3X1_129 gnd vdd FILL
XFILL_4_INVX1_10 gnd vdd FILL
XFILL_4_INVX1_21 gnd vdd FILL
XFILL_47_DFFSR_186 gnd vdd FILL
XFILL_12_NAND3X1_51 gnd vdd FILL
XFILL_12_NAND3X1_62 gnd vdd FILL
XFILL_47_DFFSR_197 gnd vdd FILL
XFILL_4_INVX1_32 gnd vdd FILL
XFILL_4_INVX1_43 gnd vdd FILL
XFILL_12_NAND3X1_73 gnd vdd FILL
XFILL_12_NAND3X1_84 gnd vdd FILL
XFILL_5_AND2X2_2 gnd vdd FILL
XFILL_12_NAND3X1_95 gnd vdd FILL
XFILL_4_INVX1_54 gnd vdd FILL
XFILL_3_BUFX2_1 gnd vdd FILL
XFILL_4_INVX1_65 gnd vdd FILL
XFILL_32_CLKBUF1_40 gnd vdd FILL
XFILL_4_INVX1_76 gnd vdd FILL
XFILL_13_AOI22X1_4 gnd vdd FILL
XFILL_4_INVX1_87 gnd vdd FILL
XFILL_4_INVX1_98 gnd vdd FILL
XFILL_11_MUX2X1_8 gnd vdd FILL
XFILL_23_MUX2X1_107 gnd vdd FILL
XFILL_23_MUX2X1_118 gnd vdd FILL
XFILL_23_MUX2X1_129 gnd vdd FILL
XFILL_17_AOI22X1_3 gnd vdd FILL
XFILL_2_BUFX4_30 gnd vdd FILL
XFILL_29_DFFSR_109 gnd vdd FILL
XFILL_2_BUFX4_41 gnd vdd FILL
XFILL_19_DFFSR_12 gnd vdd FILL
XFILL_2_BUFX4_52 gnd vdd FILL
XFILL_19_DFFSR_23 gnd vdd FILL
XFILL_2_BUFX4_63 gnd vdd FILL
XFILL_19_DFFSR_34 gnd vdd FILL
XFILL_2_BUFX4_74 gnd vdd FILL
XFILL_2_BUFX4_85 gnd vdd FILL
XFILL_19_DFFSR_45 gnd vdd FILL
XFILL_19_DFFSR_56 gnd vdd FILL
XFILL_3_OAI22X1_14 gnd vdd FILL
XFILL_2_BUFX4_96 gnd vdd FILL
XFILL_19_DFFSR_67 gnd vdd FILL
XFILL_3_OAI22X1_25 gnd vdd FILL
XFILL_19_DFFSR_78 gnd vdd FILL
XFILL_3_OAI22X1_36 gnd vdd FILL
XFILL_19_DFFSR_89 gnd vdd FILL
XFILL_3_OAI22X1_47 gnd vdd FILL
XFILL_7_OAI21X1_16 gnd vdd FILL
XFILL_59_DFFSR_11 gnd vdd FILL
XFILL_59_DFFSR_22 gnd vdd FILL
XFILL_19_2_1 gnd vdd FILL
XFILL_7_OAI21X1_27 gnd vdd FILL
XFILL_59_DFFSR_33 gnd vdd FILL
XFILL_7_OAI21X1_38 gnd vdd FILL
XFILL_7_OAI21X1_49 gnd vdd FILL
XFILL_59_DFFSR_44 gnd vdd FILL
XFILL_59_DFFSR_55 gnd vdd FILL
XFILL_59_DFFSR_66 gnd vdd FILL
XFILL_20_MUX2X1_6 gnd vdd FILL
XFILL_59_DFFSR_77 gnd vdd FILL
XFILL_62_5_2 gnd vdd FILL
XFILL_59_DFFSR_88 gnd vdd FILL
XFILL_59_DFFSR_99 gnd vdd FILL
XFILL_61_0_1 gnd vdd FILL
XFILL_10_DFFSR_110 gnd vdd FILL
XFILL_2_NAND3X1_90 gnd vdd FILL
XFILL_27_DFFSR_3 gnd vdd FILL
XFILL_0_NOR2X1_205 gnd vdd FILL
XFILL_10_DFFSR_121 gnd vdd FILL
XFILL_84_DFFSR_4 gnd vdd FILL
XFILL_4_NOR2X1_9 gnd vdd FILL
XFILL_10_DFFSR_132 gnd vdd FILL
XFILL_6_NAND2X1_70 gnd vdd FILL
XFILL_10_DFFSR_143 gnd vdd FILL
XFILL_6_NAND2X1_81 gnd vdd FILL
XFILL_28_DFFSR_10 gnd vdd FILL
XFILL_10_DFFSR_154 gnd vdd FILL
XFILL_28_DFFSR_21 gnd vdd FILL
XFILL_6_NAND2X1_92 gnd vdd FILL
XFILL_10_DFFSR_165 gnd vdd FILL
XFILL_28_DFFSR_32 gnd vdd FILL
XFILL_28_DFFSR_43 gnd vdd FILL
XFILL_3_INVX2_1 gnd vdd FILL
XFILL_12_4 gnd vdd FILL
XFILL_10_DFFSR_176 gnd vdd FILL
XFILL_10_DFFSR_187 gnd vdd FILL
XFILL_28_DFFSR_54 gnd vdd FILL
XFILL_14_CLKBUF1_12 gnd vdd FILL
XFILL_10_DFFSR_198 gnd vdd FILL
XFILL_28_DFFSR_65 gnd vdd FILL
XFILL_28_DFFSR_76 gnd vdd FILL
XFILL_14_DFFSR_120 gnd vdd FILL
XFILL_14_CLKBUF1_23 gnd vdd FILL
XFILL_28_DFFSR_87 gnd vdd FILL
XFILL_79_DFFSR_209 gnd vdd FILL
XFILL_14_DFFSR_131 gnd vdd FILL
XFILL_28_DFFSR_98 gnd vdd FILL
XFILL_14_CLKBUF1_34 gnd vdd FILL
XFILL_14_DFFSR_142 gnd vdd FILL
XFILL_14_DFFSR_153 gnd vdd FILL
XFILL_68_DFFSR_20 gnd vdd FILL
XFILL_68_DFFSR_31 gnd vdd FILL
XFILL_14_DFFSR_164 gnd vdd FILL
XFILL_68_DFFSR_42 gnd vdd FILL
XFILL_3_MUX2X1_7 gnd vdd FILL
XFILL_3_CLKBUF1_7 gnd vdd FILL
XFILL_14_DFFSR_175 gnd vdd FILL
XFILL_68_DFFSR_53 gnd vdd FILL
XFILL_14_DFFSR_186 gnd vdd FILL
XFILL_14_DFFSR_197 gnd vdd FILL
XFILL_68_DFFSR_64 gnd vdd FILL
XFILL_68_DFFSR_75 gnd vdd FILL
XFILL_18_DFFSR_130 gnd vdd FILL
XFILL_11_DFFSR_9 gnd vdd FILL
XFILL_68_DFFSR_86 gnd vdd FILL
XFILL_68_DFFSR_97 gnd vdd FILL
XFILL_18_DFFSR_141 gnd vdd FILL
XFILL_18_DFFSR_152 gnd vdd FILL
XFILL_18_DFFSR_163 gnd vdd FILL
XFILL_18_DFFSR_174 gnd vdd FILL
XFILL_10_NOR3X1_10 gnd vdd FILL
XFILL_49_DFFSR_7 gnd vdd FILL
XFILL_7_CLKBUF1_6 gnd vdd FILL
XFILL_18_DFFSR_185 gnd vdd FILL
XFILL_10_NOR3X1_21 gnd vdd FILL
XFILL_10_NOR3X1_32 gnd vdd FILL
XFILL_18_DFFSR_196 gnd vdd FILL
XFILL_37_DFFSR_30 gnd vdd FILL
XFILL_10_NOR3X1_43 gnd vdd FILL
XFILL_37_DFFSR_41 gnd vdd FILL
XFILL_60_DFFSR_210 gnd vdd FILL
XFILL_37_DFFSR_52 gnd vdd FILL
XFILL_37_DFFSR_63 gnd vdd FILL
XFILL_60_DFFSR_221 gnd vdd FILL
XFILL_3_BUFX4_101 gnd vdd FILL
XFILL_60_DFFSR_232 gnd vdd FILL
XFILL_37_DFFSR_74 gnd vdd FILL
XFILL_60_DFFSR_243 gnd vdd FILL
XFILL_37_DFFSR_85 gnd vdd FILL
XFILL_60_DFFSR_254 gnd vdd FILL
XFILL_37_DFFSR_96 gnd vdd FILL
XFILL_60_DFFSR_265 gnd vdd FILL
XFILL_14_NOR3X1_20 gnd vdd FILL
XFILL_14_NOR3X1_31 gnd vdd FILL
XFILL_14_NOR3X1_42 gnd vdd FILL
XFILL_77_DFFSR_40 gnd vdd FILL
XFILL_77_DFFSR_51 gnd vdd FILL
XFILL_77_DFFSR_62 gnd vdd FILL
XFILL_64_DFFSR_220 gnd vdd FILL
XFILL_77_DFFSR_73 gnd vdd FILL
XFILL_64_DFFSR_231 gnd vdd FILL
XFILL_7_BUFX4_100 gnd vdd FILL
XFILL_64_DFFSR_242 gnd vdd FILL
XFILL_77_DFFSR_84 gnd vdd FILL
XFILL_77_DFFSR_95 gnd vdd FILL
XFILL_64_DFFSR_253 gnd vdd FILL
XFILL_64_DFFSR_264 gnd vdd FILL
XFILL_64_DFFSR_275 gnd vdd FILL
XFILL_18_NOR3X1_30 gnd vdd FILL
XFILL_4_CLKBUF1_40 gnd vdd FILL
XFILL_18_NOR3X1_41 gnd vdd FILL
XFILL_12_MUX2X1_103 gnd vdd FILL
XFILL_18_NOR3X1_52 gnd vdd FILL
XFILL_12_MUX2X1_114 gnd vdd FILL
XFILL_53_5_2 gnd vdd FILL
XFILL_12_MUX2X1_125 gnd vdd FILL
XFILL_0_INVX1_80 gnd vdd FILL
XFILL_0_INVX1_91 gnd vdd FILL
XFILL_68_DFFSR_230 gnd vdd FILL
XFILL_17_NOR3X1_3 gnd vdd FILL
XFILL_68_DFFSR_241 gnd vdd FILL
XFILL_12_MUX2X1_136 gnd vdd FILL
XFILL_52_0_1 gnd vdd FILL
XFILL_68_DFFSR_252 gnd vdd FILL
XFILL_12_MUX2X1_147 gnd vdd FILL
XFILL_12_MUX2X1_158 gnd vdd FILL
XFILL_46_DFFSR_50 gnd vdd FILL
XFILL_12_MUX2X1_169 gnd vdd FILL
XFILL_46_DFFSR_61 gnd vdd FILL
XFILL_68_DFFSR_263 gnd vdd FILL
XFILL_68_DFFSR_274 gnd vdd FILL
XFILL_23_CLKBUF1_4 gnd vdd FILL
XFILL_46_DFFSR_72 gnd vdd FILL
XFILL_46_DFFSR_83 gnd vdd FILL
XFILL_1_NOR2X1_14 gnd vdd FILL
XFILL_1_NOR2X1_25 gnd vdd FILL
XFILL_46_DFFSR_94 gnd vdd FILL
XFILL_13_OAI21X1_30 gnd vdd FILL
XFILL_1_NOR2X1_36 gnd vdd FILL
XFILL_1_NOR2X1_47 gnd vdd FILL
XFILL_13_OAI21X1_41 gnd vdd FILL
XFILL_1_NOR2X1_58 gnd vdd FILL
XFILL_1_NOR2X1_69 gnd vdd FILL
XFILL_27_CLKBUF1_3 gnd vdd FILL
XFILL_86_DFFSR_60 gnd vdd FILL
XFILL_2_NOR2X1_180 gnd vdd FILL
XFILL_86_DFFSR_71 gnd vdd FILL
XFILL_86_DFFSR_82 gnd vdd FILL
XFILL_86_DFFSR_93 gnd vdd FILL
XFILL_2_NOR2X1_191 gnd vdd FILL
XFILL_5_NOR2X1_13 gnd vdd FILL
XFILL_5_NOR2X1_24 gnd vdd FILL
XFILL_46_DFFSR_209 gnd vdd FILL
XFILL_15_DFFSR_60 gnd vdd FILL
XFILL_5_NOR2X1_35 gnd vdd FILL
XFILL_15_DFFSR_71 gnd vdd FILL
XFILL_15_DFFSR_82 gnd vdd FILL
XFILL_5_NOR2X1_46 gnd vdd FILL
XFILL_15_DFFSR_93 gnd vdd FILL
XFILL_5_NOR2X1_57 gnd vdd FILL
XFILL_5_NOR2X1_68 gnd vdd FILL
XFILL_5_NOR2X1_79 gnd vdd FILL
XFILL_26_NOR3X1_1 gnd vdd FILL
XFILL_73_DFFSR_109 gnd vdd FILL
XFILL_9_NOR2X1_12 gnd vdd FILL
XFILL_9_NOR2X1_23 gnd vdd FILL
XFILL_9_NOR2X1_34 gnd vdd FILL
XFILL_55_DFFSR_70 gnd vdd FILL
XFILL_55_DFFSR_81 gnd vdd FILL
XFILL_9_NOR2X1_45 gnd vdd FILL
XFILL_9_NOR2X1_56 gnd vdd FILL
XFILL_55_DFFSR_92 gnd vdd FILL
XFILL_13_OAI22X1_7 gnd vdd FILL
XFILL_9_NOR2X1_67 gnd vdd FILL
XFILL_9_NOR2X1_78 gnd vdd FILL
XFILL_9_NOR2X1_89 gnd vdd FILL
XFILL_0_NOR2X1_2 gnd vdd FILL
XFILL_2_MUX2X1_120 gnd vdd FILL
XFILL_77_DFFSR_108 gnd vdd FILL
XFILL_77_DFFSR_119 gnd vdd FILL
XFILL_2_MUX2X1_131 gnd vdd FILL
XFILL_2_MUX2X1_142 gnd vdd FILL
XFILL_2_MUX2X1_153 gnd vdd FILL
XFILL_17_OAI22X1_6 gnd vdd FILL
XFILL_2_MUX2X1_164 gnd vdd FILL
XFILL_15_NAND3X1_17 gnd vdd FILL
XFILL_2_MUX2X1_175 gnd vdd FILL
XFILL_15_NAND3X1_28 gnd vdd FILL
XFILL_2_MUX2X1_186 gnd vdd FILL
XFILL_15_NAND3X1_39 gnd vdd FILL
XFILL_24_DFFSR_80 gnd vdd FILL
XFILL_24_DFFSR_91 gnd vdd FILL
XFILL_9_NOR3X1_2 gnd vdd FILL
XFILL_35_CLKBUF1_17 gnd vdd FILL
XFILL_35_CLKBUF1_28 gnd vdd FILL
XFILL_31_DFFSR_220 gnd vdd FILL
XFILL_7_BUFX2_2 gnd vdd FILL
XFILL_31_DFFSR_231 gnd vdd FILL
XFILL_35_CLKBUF1_39 gnd vdd FILL
XFILL_31_DFFSR_242 gnd vdd FILL
XFILL_31_DFFSR_253 gnd vdd FILL
XFILL_44_5_2 gnd vdd FILL
XFILL_31_DFFSR_264 gnd vdd FILL
XFILL_31_DFFSR_275 gnd vdd FILL
XFILL_64_DFFSR_90 gnd vdd FILL
XFILL_43_0_1 gnd vdd FILL
XFILL_35_DFFSR_230 gnd vdd FILL
XFILL_35_DFFSR_241 gnd vdd FILL
XFILL_66_DFFSR_1 gnd vdd FILL
XFILL_35_DFFSR_252 gnd vdd FILL
XFILL_1_MUX2X1_10 gnd vdd FILL
XFILL_35_DFFSR_263 gnd vdd FILL
XFILL_35_DFFSR_274 gnd vdd FILL
XFILL_1_MUX2X1_21 gnd vdd FILL
XFILL_7_DFFSR_70 gnd vdd FILL
XFILL_1_MUX2X1_32 gnd vdd FILL
XFILL_7_DFFSR_81 gnd vdd FILL
XFILL_7_DFFSR_92 gnd vdd FILL
XFILL_1_MUX2X1_43 gnd vdd FILL
XFILL_1_MUX2X1_54 gnd vdd FILL
XFILL_62_DFFSR_130 gnd vdd FILL
XFILL_1_MUX2X1_65 gnd vdd FILL
XFILL_1_MUX2X1_76 gnd vdd FILL
XFILL_39_DFFSR_240 gnd vdd FILL
XFILL_62_DFFSR_141 gnd vdd FILL
XFILL_62_DFFSR_152 gnd vdd FILL
XFILL_39_DFFSR_251 gnd vdd FILL
XFILL_1_MUX2X1_87 gnd vdd FILL
XFILL_14_NAND3X1_108 gnd vdd FILL
XFILL_62_DFFSR_163 gnd vdd FILL
XFILL_62_DFFSR_174 gnd vdd FILL
XFILL_39_DFFSR_262 gnd vdd FILL
XFILL_14_NAND3X1_119 gnd vdd FILL
XFILL_1_MUX2X1_98 gnd vdd FILL
XFILL_39_DFFSR_273 gnd vdd FILL
XFILL_5_MUX2X1_20 gnd vdd FILL
XFILL_5_MUX2X1_31 gnd vdd FILL
XFILL_62_DFFSR_185 gnd vdd FILL
XFILL_62_DFFSR_196 gnd vdd FILL
XFILL_5_NAND3X1_12 gnd vdd FILL
XFILL_5_MUX2X1_42 gnd vdd FILL
XFILL_13_DFFSR_209 gnd vdd FILL
XFILL_5_MUX2X1_53 gnd vdd FILL
XFILL_10_NAND3X1_9 gnd vdd FILL
XFILL_5_MUX2X1_64 gnd vdd FILL
XFILL_5_NAND3X1_23 gnd vdd FILL
XFILL_66_DFFSR_140 gnd vdd FILL
XFILL_5_MUX2X1_75 gnd vdd FILL
XFILL_5_NAND3X1_34 gnd vdd FILL
XFILL_66_DFFSR_151 gnd vdd FILL
XFILL_5_NAND3X1_45 gnd vdd FILL
XFILL_66_DFFSR_162 gnd vdd FILL
XFILL_5_MUX2X1_86 gnd vdd FILL
XFILL_5_NAND3X1_56 gnd vdd FILL
XFILL_5_MUX2X1_97 gnd vdd FILL
XFILL_9_NAND2X1_14 gnd vdd FILL
XFILL_66_DFFSR_173 gnd vdd FILL
XFILL_5_NAND3X1_67 gnd vdd FILL
XFILL_50_DFFSR_7 gnd vdd FILL
XFILL_66_DFFSR_184 gnd vdd FILL
XFILL_9_NAND2X1_25 gnd vdd FILL
XFILL_9_MUX2X1_30 gnd vdd FILL
XFILL_5_NAND3X1_78 gnd vdd FILL
XFILL_9_NAND2X1_36 gnd vdd FILL
XFILL_40_DFFSR_109 gnd vdd FILL
XFILL_5_NAND3X1_89 gnd vdd FILL
XFILL_66_DFFSR_195 gnd vdd FILL
XFILL_9_MUX2X1_41 gnd vdd FILL
XFILL_9_NAND2X1_47 gnd vdd FILL
XFILL_17_DFFSR_208 gnd vdd FILL
XFILL_14_NAND3X1_8 gnd vdd FILL
XFILL_17_DFFSR_219 gnd vdd FILL
XFILL_9_MUX2X1_52 gnd vdd FILL
XFILL_9_NAND2X1_58 gnd vdd FILL
XFILL_9_NAND2X1_69 gnd vdd FILL
XFILL_9_MUX2X1_63 gnd vdd FILL
XFILL_9_MUX2X1_74 gnd vdd FILL
XFILL_9_MUX2X1_85 gnd vdd FILL
XFILL_7_INVX2_2 gnd vdd FILL
XFILL_9_MUX2X1_96 gnd vdd FILL
XFILL_44_DFFSR_108 gnd vdd FILL
XBUFX4_20 BUFX4_3/Y gnd DFFSR_78/R vdd BUFX4
XFILL_44_DFFSR_119 gnd vdd FILL
XFILL_67_5 gnd vdd FILL
XBUFX4_31 BUFX4_44/A gnd DFFSR_79/R vdd BUFX4
XBUFX4_42 BUFX4_44/A gnd DFFSR_48/R vdd BUFX4
XBUFX4_53 BUFX4_54/A gnd DFFSR_9/R vdd BUFX4
XFILL_12_AOI21X1_19 gnd vdd FILL
XBUFX4_64 INVX8_1/Y gnd BUFX4_64/Y vdd BUFX4
XBUFX4_75 INVX8_2/Y gnd BUFX4_75/Y vdd BUFX4
XBUFX4_86 INVX8_4/Y gnd BUFX4_86/Y vdd BUFX4
XBUFX4_97 INVX8_3/Y gnd BUFX4_97/Y vdd BUFX4
XFILL_48_DFFSR_107 gnd vdd FILL
XFILL_48_DFFSR_118 gnd vdd FILL
XFILL_3_BUFX4_19 gnd vdd FILL
XFILL_48_DFFSR_129 gnd vdd FILL
XFILL_35_5_2 gnd vdd FILL
XFILL_21_MUX2X1_40 gnd vdd FILL
XFILL_21_MUX2X1_51 gnd vdd FILL
XFILL_21_MUX2X1_62 gnd vdd FILL
XFILL_21_MUX2X1_73 gnd vdd FILL
XFILL_34_0_1 gnd vdd FILL
XFILL_21_MUX2X1_84 gnd vdd FILL
XFILL_21_MUX2X1_95 gnd vdd FILL
XFILL_10_1 gnd vdd FILL
XFILL_24_CLKBUF1_13 gnd vdd FILL
XFILL_24_CLKBUF1_24 gnd vdd FILL
XFILL_24_CLKBUF1_35 gnd vdd FILL
XFILL_0_NAND3X1_109 gnd vdd FILL
XFILL_7_CLKBUF1_17 gnd vdd FILL
XFILL_7_CLKBUF1_28 gnd vdd FILL
XFILL_10_AND2X2_7 gnd vdd FILL
XFILL_7_CLKBUF1_39 gnd vdd FILL
XFILL_2_AOI21X1_14 gnd vdd FILL
XFILL_2_AOI21X1_25 gnd vdd FILL
XFILL_33_DFFSR_140 gnd vdd FILL
XFILL_2_AOI21X1_36 gnd vdd FILL
XFILL_33_DFFSR_151 gnd vdd FILL
XFILL_33_DFFSR_162 gnd vdd FILL
XFILL_2_AOI21X1_47 gnd vdd FILL
XFILL_33_DFFSR_173 gnd vdd FILL
XFILL_12_OAI22X1_16 gnd vdd FILL
XFILL_2_AOI21X1_58 gnd vdd FILL
XFILL_2_AOI21X1_69 gnd vdd FILL
XFILL_33_DFFSR_184 gnd vdd FILL
XFILL_12_OAI22X1_27 gnd vdd FILL
XFILL_33_DFFSR_195 gnd vdd FILL
XFILL_12_OAI22X1_38 gnd vdd FILL
XFILL_5_NOR2X1_102 gnd vdd FILL
XFILL_12_OAI22X1_49 gnd vdd FILL
XFILL_5_NOR2X1_113 gnd vdd FILL
XFILL_5_NOR2X1_124 gnd vdd FILL
XFILL_37_DFFSR_150 gnd vdd FILL
XFILL_5_NOR2X1_135 gnd vdd FILL
XFILL_37_DFFSR_161 gnd vdd FILL
XFILL_5_NOR2X1_146 gnd vdd FILL
XFILL_5_NOR2X1_157 gnd vdd FILL
XFILL_37_DFFSR_172 gnd vdd FILL
XFILL_37_DFFSR_183 gnd vdd FILL
XFILL_5_NOR2X1_168 gnd vdd FILL
XFILL_5_NOR2X1_179 gnd vdd FILL
XFILL_11_DFFSR_108 gnd vdd FILL
XFILL_37_DFFSR_194 gnd vdd FILL
XFILL_11_NAND3X1_70 gnd vdd FILL
XFILL_11_NAND3X1_81 gnd vdd FILL
XFILL_11_DFFSR_119 gnd vdd FILL
XFILL_11_NAND3X1_92 gnd vdd FILL
XFILL_38_DFFSR_19 gnd vdd FILL
XFILL_1_5_2 gnd vdd FILL
XFILL_26_5_2 gnd vdd FILL
XFILL_15_DFFSR_107 gnd vdd FILL
XFILL_15_DFFSR_118 gnd vdd FILL
XFILL_25_0_1 gnd vdd FILL
XFILL_22_MUX2X1_104 gnd vdd FILL
XFILL_0_0_1 gnd vdd FILL
XFILL_22_MUX2X1_115 gnd vdd FILL
XFILL_15_DFFSR_129 gnd vdd FILL
XFILL_22_MUX2X1_126 gnd vdd FILL
XFILL_10_AOI21X1_3 gnd vdd FILL
XFILL_78_DFFSR_18 gnd vdd FILL
XFILL_78_DFFSR_29 gnd vdd FILL
XFILL_22_MUX2X1_137 gnd vdd FILL
XFILL_83_DFFSR_240 gnd vdd FILL
XFILL_22_MUX2X1_148 gnd vdd FILL
XFILL_22_MUX2X1_159 gnd vdd FILL
XFILL_83_DFFSR_251 gnd vdd FILL
XFILL_83_DFFSR_262 gnd vdd FILL
XFILL_19_DFFSR_106 gnd vdd FILL
XFILL_83_DFFSR_273 gnd vdd FILL
XFILL_5_MUX2X1_108 gnd vdd FILL
XFILL_5_MUX2X1_119 gnd vdd FILL
XFILL_19_DFFSR_117 gnd vdd FILL
XFILL_19_DFFSR_128 gnd vdd FILL
XFILL_1_INVX1_14 gnd vdd FILL
XFILL_1_INVX1_25 gnd vdd FILL
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XFILL_1_INVX1_36 gnd vdd FILL
XFILL_19_DFFSR_139 gnd vdd FILL
XFILL_14_AOI21X1_2 gnd vdd FILL
XFILL_2_OAI22X1_11 gnd vdd FILL
XFILL_1_INVX1_47 gnd vdd FILL
XFILL_2_OAI22X1_22 gnd vdd FILL
XFILL_2_AND2X2_6 gnd vdd FILL
XFILL_1_INVX1_58 gnd vdd FILL
XFILL_2_OAI22X1_33 gnd vdd FILL
XFILL_87_DFFSR_250 gnd vdd FILL
XFILL_2_OAI22X1_44 gnd vdd FILL
XFILL_1_INVX1_69 gnd vdd FILL
XFILL_47_DFFSR_17 gnd vdd FILL
XFILL_11_NOR3X1_19 gnd vdd FILL
XFILL_87_DFFSR_261 gnd vdd FILL
XFILL_6_OAI21X1_13 gnd vdd FILL
XFILL_87_DFFSR_272 gnd vdd FILL
XFILL_6_OAI21X1_24 gnd vdd FILL
XFILL_47_DFFSR_28 gnd vdd FILL
XFILL_47_DFFSR_39 gnd vdd FILL
XFILL_61_DFFSR_208 gnd vdd FILL
XFILL_6_OAI21X1_35 gnd vdd FILL
XFILL_61_DFFSR_219 gnd vdd FILL
XFILL_6_OAI21X1_46 gnd vdd FILL
XFILL_15_NOR3X1_18 gnd vdd FILL
XFILL_87_DFFSR_16 gnd vdd FILL
XFILL_87_DFFSR_27 gnd vdd FILL
XFILL_15_NOR3X1_29 gnd vdd FILL
XFILL_32_DFFSR_4 gnd vdd FILL
XFILL_87_DFFSR_38 gnd vdd FILL
XFILL_65_DFFSR_207 gnd vdd FILL
XFILL_87_DFFSR_49 gnd vdd FILL
XFILL_16_DFFSR_16 gnd vdd FILL
XFILL_65_DFFSR_218 gnd vdd FILL
XFILL_9_6_2 gnd vdd FILL
XFILL_16_DFFSR_27 gnd vdd FILL
XFILL_65_DFFSR_229 gnd vdd FILL
XFILL_16_DFFSR_38 gnd vdd FILL
XFILL_8_1_1 gnd vdd FILL
XFILL_16_DFFSR_49 gnd vdd FILL
XFILL_19_NOR3X1_17 gnd vdd FILL
XFILL_19_NOR3X1_28 gnd vdd FILL
XFILL_19_NOR3X1_39 gnd vdd FILL
XFILL_13_CLKBUF1_20 gnd vdd FILL
XFILL_69_DFFSR_206 gnd vdd FILL
XFILL_13_CLKBUF1_31 gnd vdd FILL
XFILL_69_DFFSR_217 gnd vdd FILL
XFILL_56_DFFSR_15 gnd vdd FILL
XFILL_56_DFFSR_26 gnd vdd FILL
XFILL_13_CLKBUF1_42 gnd vdd FILL
XFILL_69_DFFSR_228 gnd vdd FILL
XFILL_56_DFFSR_37 gnd vdd FILL
XFILL_69_DFFSR_239 gnd vdd FILL
XFILL_56_DFFSR_48 gnd vdd FILL
XFILL_56_DFFSR_59 gnd vdd FILL
XFILL_17_5_2 gnd vdd FILL
XFILL_54_DFFSR_8 gnd vdd FILL
XFILL_16_0_1 gnd vdd FILL
XFILL_25_DFFSR_14 gnd vdd FILL
XFILL_25_DFFSR_25 gnd vdd FILL
XFILL_11_NOR2X1_160 gnd vdd FILL
XFILL_25_DFFSR_36 gnd vdd FILL
XFILL_25_DFFSR_47 gnd vdd FILL
XFILL_11_NOR2X1_171 gnd vdd FILL
XFILL_25_DFFSR_58 gnd vdd FILL
XFILL_11_NOR2X1_182 gnd vdd FILL
XFILL_11_NOR2X1_193 gnd vdd FILL
XFILL_25_DFFSR_69 gnd vdd FILL
XFILL_50_DFFSR_240 gnd vdd FILL
XFILL_65_DFFSR_13 gnd vdd FILL
XFILL_50_DFFSR_251 gnd vdd FILL
XFILL_65_DFFSR_24 gnd vdd FILL
XFILL_50_DFFSR_262 gnd vdd FILL
XFILL_65_DFFSR_35 gnd vdd FILL
XFILL_50_DFFSR_273 gnd vdd FILL
XFILL_65_DFFSR_46 gnd vdd FILL
XFILL_65_DFFSR_57 gnd vdd FILL
XFILL_65_DFFSR_68 gnd vdd FILL
XFILL_65_DFFSR_79 gnd vdd FILL
XFILL_54_DFFSR_250 gnd vdd FILL
XFILL_15_NAND3X1_109 gnd vdd FILL
XFILL_54_DFFSR_261 gnd vdd FILL
XFILL_54_DFFSR_272 gnd vdd FILL
XFILL_8_DFFSR_15 gnd vdd FILL
XFILL_8_DFFSR_26 gnd vdd FILL
XFILL_11_MUX2X1_100 gnd vdd FILL
XFILL_34_DFFSR_12 gnd vdd FILL
XFILL_8_DFFSR_37 gnd vdd FILL
XFILL_11_MUX2X1_111 gnd vdd FILL
XFILL_8_DFFSR_48 gnd vdd FILL
XFILL_11_MUX2X1_122 gnd vdd FILL
XFILL_34_DFFSR_23 gnd vdd FILL
XFILL_34_DFFSR_34 gnd vdd FILL
XFILL_8_DFFSR_59 gnd vdd FILL
XFILL_34_DFFSR_45 gnd vdd FILL
XFILL_11_MUX2X1_133 gnd vdd FILL
XFILL_11_MUX2X1_144 gnd vdd FILL
XFILL_34_DFFSR_56 gnd vdd FILL
XFILL_81_DFFSR_150 gnd vdd FILL
XFILL_81_DFFSR_161 gnd vdd FILL
XFILL_11_MUX2X1_155 gnd vdd FILL
XFILL_34_DFFSR_67 gnd vdd FILL
XFILL_13_CLKBUF1_1 gnd vdd FILL
XFILL_81_DFFSR_172 gnd vdd FILL
XFILL_58_DFFSR_260 gnd vdd FILL
XFILL_11_MUX2X1_166 gnd vdd FILL
XFILL_58_DFFSR_271 gnd vdd FILL
XFILL_34_DFFSR_78 gnd vdd FILL
XFILL_11_MUX2X1_177 gnd vdd FILL
XFILL_34_DFFSR_89 gnd vdd FILL
XFILL_81_DFFSR_183 gnd vdd FILL
XFILL_74_DFFSR_11 gnd vdd FILL
XFILL_11_MUX2X1_188 gnd vdd FILL
XFILL_81_DFFSR_194 gnd vdd FILL
XFILL_32_DFFSR_207 gnd vdd FILL
XFILL_1_DFFSR_220 gnd vdd FILL
XFILL_74_DFFSR_22 gnd vdd FILL
XFILL_32_DFFSR_218 gnd vdd FILL
XFILL_1_DFFSR_231 gnd vdd FILL
XFILL_1_DFFSR_242 gnd vdd FILL
XFILL_32_DFFSR_229 gnd vdd FILL
XFILL_74_DFFSR_33 gnd vdd FILL
XFILL_17_MUX2X1_1 gnd vdd FILL
XFILL_74_DFFSR_44 gnd vdd FILL
XFILL_74_DFFSR_55 gnd vdd FILL
XFILL_1_DFFSR_253 gnd vdd FILL
XFILL_85_DFFSR_160 gnd vdd FILL
XFILL_74_DFFSR_66 gnd vdd FILL
XFILL_1_DFFSR_264 gnd vdd FILL
XFILL_1_DFFSR_275 gnd vdd FILL
XFILL_74_DFFSR_77 gnd vdd FILL
XFILL_85_DFFSR_171 gnd vdd FILL
XFILL_65_2 gnd vdd FILL
XFILL_85_DFFSR_182 gnd vdd FILL
XFILL_74_DFFSR_88 gnd vdd FILL
XFILL_74_DFFSR_99 gnd vdd FILL
XFILL_85_DFFSR_193 gnd vdd FILL
XFILL_36_DFFSR_206 gnd vdd FILL
XFILL_36_DFFSR_217 gnd vdd FILL
XFILL_5_DFFSR_230 gnd vdd FILL
XFILL_58_1 gnd vdd FILL
XFILL_5_DFFSR_241 gnd vdd FILL
XFILL_36_DFFSR_228 gnd vdd FILL
XFILL_36_DFFSR_239 gnd vdd FILL
XFILL_5_DFFSR_252 gnd vdd FILL
XFILL_43_DFFSR_10 gnd vdd FILL
XFILL_43_DFFSR_21 gnd vdd FILL
XFILL_5_DFFSR_263 gnd vdd FILL
XFILL_5_DFFSR_274 gnd vdd FILL
XFILL_43_DFFSR_32 gnd vdd FILL
XFILL_2_MUX2X1_19 gnd vdd FILL
XFILL_14_NOR3X1_7 gnd vdd FILL
XFILL_43_DFFSR_43 gnd vdd FILL
XFILL_63_DFFSR_106 gnd vdd FILL
XFILL_43_DFFSR_54 gnd vdd FILL
XFILL_43_DFFSR_65 gnd vdd FILL
XFILL_63_DFFSR_117 gnd vdd FILL
XFILL_43_DFFSR_76 gnd vdd FILL
XFILL_43_DFFSR_87 gnd vdd FILL
XFILL_9_DFFSR_240 gnd vdd FILL
XFILL_63_DFFSR_128 gnd vdd FILL
XFILL_9_DFFSR_251 gnd vdd FILL
XFILL_63_DFFSR_139 gnd vdd FILL
XFILL_43_DFFSR_98 gnd vdd FILL
XFILL_10_NAND3X1_105 gnd vdd FILL
XFILL_10_NAND3X1_116 gnd vdd FILL
XFILL_9_DFFSR_262 gnd vdd FILL
XFILL_83_DFFSR_20 gnd vdd FILL
XFILL_9_DFFSR_273 gnd vdd FILL
XFILL_83_DFFSR_31 gnd vdd FILL
XFILL_10_NAND3X1_127 gnd vdd FILL
XFILL_6_MUX2X1_18 gnd vdd FILL
XFILL_83_DFFSR_42 gnd vdd FILL
XFILL_50_3_2 gnd vdd FILL
XFILL_6_MUX2X1_29 gnd vdd FILL
XFILL_67_DFFSR_105 gnd vdd FILL
XFILL_83_DFFSR_53 gnd vdd FILL
XFILL_12_DFFSR_20 gnd vdd FILL
XFILL_67_DFFSR_116 gnd vdd FILL
XFILL_83_DFFSR_64 gnd vdd FILL
XFILL_67_DFFSR_127 gnd vdd FILL
XFILL_12_DFFSR_31 gnd vdd FILL
XFILL_83_DFFSR_75 gnd vdd FILL
XFILL_83_DFFSR_86 gnd vdd FILL
XFILL_1_MUX2X1_150 gnd vdd FILL
XFILL_12_DFFSR_42 gnd vdd FILL
XFILL_67_DFFSR_138 gnd vdd FILL
XFILL_83_DFFSR_97 gnd vdd FILL
XFILL_1_MUX2X1_161 gnd vdd FILL
XFILL_67_DFFSR_149 gnd vdd FILL
XFILL_10_OAI21X1_6 gnd vdd FILL
XFILL_14_NAND3X1_14 gnd vdd FILL
XFILL_12_DFFSR_53 gnd vdd FILL
XFILL_14_NAND3X1_25 gnd vdd FILL
XFILL_1_MUX2X1_172 gnd vdd FILL
XFILL_12_DFFSR_64 gnd vdd FILL
XFILL_12_DFFSR_75 gnd vdd FILL
XFILL_14_NAND3X1_36 gnd vdd FILL
XFILL_1_MUX2X1_183 gnd vdd FILL
XFILL_12_DFFSR_86 gnd vdd FILL
XFILL_1_MUX2X1_194 gnd vdd FILL
XFILL_14_NAND3X1_47 gnd vdd FILL
XFILL_12_DFFSR_97 gnd vdd FILL
XFILL_14_NAND3X1_58 gnd vdd FILL
XFILL_14_NAND3X1_69 gnd vdd FILL
XFILL_34_CLKBUF1_14 gnd vdd FILL
XFILL_34_CLKBUF1_25 gnd vdd FILL
XFILL_52_DFFSR_30 gnd vdd FILL
XFILL_34_CLKBUF1_36 gnd vdd FILL
XFILL_52_DFFSR_41 gnd vdd FILL
XFILL_23_NOR3X1_5 gnd vdd FILL
XFILL_11_NOR2X1_30 gnd vdd FILL
XFILL_2_AOI22X1_2 gnd vdd FILL
XFILL_52_DFFSR_52 gnd vdd FILL
XFILL_14_OAI21X1_5 gnd vdd FILL
XFILL_52_DFFSR_63 gnd vdd FILL
XFILL_11_NOR2X1_41 gnd vdd FILL
XFILL_11_NOR2X1_52 gnd vdd FILL
XFILL_52_DFFSR_74 gnd vdd FILL
XFILL_21_DFFSR_250 gnd vdd FILL
XFILL_52_DFFSR_85 gnd vdd FILL
XFILL_11_NOR2X1_63 gnd vdd FILL
XFILL_21_DFFSR_261 gnd vdd FILL
XFILL_21_DFFSR_272 gnd vdd FILL
XFILL_11_NOR2X1_74 gnd vdd FILL
XFILL_52_DFFSR_96 gnd vdd FILL
XFILL_11_NOR2X1_85 gnd vdd FILL
XFILL_2_INVX1_201 gnd vdd FILL
XFILL_1_DFFSR_3 gnd vdd FILL
XFILL_2_INVX1_212 gnd vdd FILL
XFILL_2_INVX1_223 gnd vdd FILL
XFILL_11_NOR2X1_96 gnd vdd FILL
XFILL_6_AOI22X1_1 gnd vdd FILL
XFILL_14_DFFSR_1 gnd vdd FILL
XFILL_71_DFFSR_2 gnd vdd FILL
XFILL_21_DFFSR_40 gnd vdd FILL
XFILL_25_DFFSR_260 gnd vdd FILL
XFILL_25_DFFSR_271 gnd vdd FILL
XFILL_21_DFFSR_51 gnd vdd FILL
XFILL_6_INVX1_200 gnd vdd FILL
XFILL_22_MUX2X1_16 gnd vdd FILL
XFILL_21_DFFSR_62 gnd vdd FILL
XFILL_22_MUX2X1_27 gnd vdd FILL
XFILL_6_INVX1_211 gnd vdd FILL
XFILL_21_DFFSR_73 gnd vdd FILL
XFILL_6_INVX1_222 gnd vdd FILL
XFILL_21_DFFSR_84 gnd vdd FILL
XFILL_22_MUX2X1_38 gnd vdd FILL
XFILL_58_4_2 gnd vdd FILL
XFILL_21_DFFSR_95 gnd vdd FILL
XFILL_22_MUX2X1_49 gnd vdd FILL
XFILL_6_NOR3X1_6 gnd vdd FILL
XFILL_52_DFFSR_160 gnd vdd FILL
XFILL_52_DFFSR_171 gnd vdd FILL
XFILL_29_DFFSR_270 gnd vdd FILL
XFILL_52_DFFSR_182 gnd vdd FILL
XFILL_61_DFFSR_50 gnd vdd FILL
XFILL_61_DFFSR_61 gnd vdd FILL
XFILL_52_DFFSR_193 gnd vdd FILL
XFILL_61_DFFSR_72 gnd vdd FILL
XFILL_61_DFFSR_83 gnd vdd FILL
XFILL_4_NAND3X1_20 gnd vdd FILL
XFILL_61_DFFSR_94 gnd vdd FILL
XFILL_4_NAND3X1_31 gnd vdd FILL
XFILL_4_NAND3X1_42 gnd vdd FILL
XFILL_4_NAND3X1_53 gnd vdd FILL
XFILL_56_DFFSR_170 gnd vdd FILL
XFILL_4_NAND3X1_64 gnd vdd FILL
XFILL_8_NAND2X1_11 gnd vdd FILL
XFILL_4_NAND3X1_75 gnd vdd FILL
XFILL_4_DFFSR_30 gnd vdd FILL
XFILL_8_NAND2X1_22 gnd vdd FILL
XFILL_56_DFFSR_181 gnd vdd FILL
XFILL_36_DFFSR_5 gnd vdd FILL
XFILL_4_DFFSR_41 gnd vdd FILL
XFILL_8_NAND2X1_33 gnd vdd FILL
XFILL_30_DFFSR_106 gnd vdd FILL
XFILL_8_NAND2X1_44 gnd vdd FILL
XFILL_4_NAND3X1_86 gnd vdd FILL
XFILL_56_DFFSR_192 gnd vdd FILL
XFILL_4_DFFSR_52 gnd vdd FILL
XFILL_4_DFFSR_63 gnd vdd FILL
XFILL_4_NAND3X1_97 gnd vdd FILL
XFILL_30_DFFSR_117 gnd vdd FILL
XFILL_8_NAND2X1_55 gnd vdd FILL
XFILL_8_NAND2X1_66 gnd vdd FILL
XFILL_4_DFFSR_74 gnd vdd FILL
XFILL_30_DFFSR_128 gnd vdd FILL
XFILL_41_3_2 gnd vdd FILL
XFILL_8_NAND2X1_77 gnd vdd FILL
XFILL_4_DFFSR_85 gnd vdd FILL
XFILL_30_DFFSR_60 gnd vdd FILL
XFILL_30_DFFSR_139 gnd vdd FILL
XFILL_4_DFFSR_96 gnd vdd FILL
XFILL_8_NAND2X1_88 gnd vdd FILL
XFILL_30_DFFSR_71 gnd vdd FILL
XFILL_30_DFFSR_82 gnd vdd FILL
XFILL_30_DFFSR_93 gnd vdd FILL
XFILL_34_DFFSR_105 gnd vdd FILL
XFILL_16_CLKBUF1_19 gnd vdd FILL
XFILL_34_DFFSR_116 gnd vdd FILL
XFILL_34_DFFSR_127 gnd vdd FILL
XFILL_11_NAND2X1_7 gnd vdd FILL
XFILL_3_DFFSR_140 gnd vdd FILL
XFILL_10_7_0 gnd vdd FILL
XFILL_34_DFFSR_138 gnd vdd FILL
XFILL_3_DFFSR_151 gnd vdd FILL
XFILL_3_DFFSR_162 gnd vdd FILL
XFILL_34_DFFSR_149 gnd vdd FILL
XFILL_11_AOI21X1_16 gnd vdd FILL
XFILL_70_DFFSR_70 gnd vdd FILL
XFILL_3_DFFSR_173 gnd vdd FILL
XFILL_11_AOI21X1_27 gnd vdd FILL
XFILL_70_DFFSR_81 gnd vdd FILL
XFILL_3_DFFSR_184 gnd vdd FILL
XFILL_70_DFFSR_92 gnd vdd FILL
XFILL_11_AOI21X1_38 gnd vdd FILL
XFILL_11_AOI21X1_49 gnd vdd FILL
XAND2X2_7 AND2X2_7/A INVX1_57/A gnd AND2X2_7/Y vdd AND2X2
XFILL_3_DFFSR_195 gnd vdd FILL
XFILL_38_DFFSR_104 gnd vdd FILL
XFILL_38_DFFSR_115 gnd vdd FILL
XFILL_38_DFFSR_126 gnd vdd FILL
XFILL_38_DFFSR_137 gnd vdd FILL
XFILL_7_DFFSR_150 gnd vdd FILL
XFILL_7_DFFSR_161 gnd vdd FILL
XFILL_38_DFFSR_148 gnd vdd FILL
XFILL_58_DFFSR_9 gnd vdd FILL
XFILL_7_DFFSR_172 gnd vdd FILL
XFILL_11_MUX2X1_70 gnd vdd FILL
XFILL_38_DFFSR_159 gnd vdd FILL
XFILL_11_MUX2X1_81 gnd vdd FILL
XFILL_7_DFFSR_183 gnd vdd FILL
XFILL_11_MUX2X1_92 gnd vdd FILL
XFILL_30_NOR3X1_17 gnd vdd FILL
XFILL_7_DFFSR_194 gnd vdd FILL
XFILL_30_NOR3X1_28 gnd vdd FILL
XFILL_30_NOR3X1_39 gnd vdd FILL
XFILL_80_DFFSR_206 gnd vdd FILL
XFILL_80_DFFSR_217 gnd vdd FILL
XFILL_80_DFFSR_228 gnd vdd FILL
XFILL_80_DFFSR_239 gnd vdd FILL
XFILL_15_MUX2X1_80 gnd vdd FILL
XFILL_15_MUX2X1_91 gnd vdd FILL
XFILL_49_4_2 gnd vdd FILL
XFILL_3_NOR3X1_40 gnd vdd FILL
XFILL_3_NOR3X1_51 gnd vdd FILL
XFILL_23_CLKBUF1_10 gnd vdd FILL
XFILL_23_CLKBUF1_21 gnd vdd FILL
XFILL_23_CLKBUF1_32 gnd vdd FILL
XFILL_84_DFFSR_205 gnd vdd FILL
XFILL_84_DFFSR_216 gnd vdd FILL
XFILL_84_DFFSR_227 gnd vdd FILL
XFILL_84_DFFSR_238 gnd vdd FILL
XFILL_84_DFFSR_249 gnd vdd FILL
XFILL_19_MUX2X1_90 gnd vdd FILL
XFILL_0_INVX1_100 gnd vdd FILL
XFILL_6_CLKBUF1_14 gnd vdd FILL
XFILL_6_CLKBUF1_25 gnd vdd FILL
XFILL_0_INVX1_111 gnd vdd FILL
XFILL_6_CLKBUF1_36 gnd vdd FILL
XFILL_7_NOR3X1_50 gnd vdd FILL
XFILL_0_INVX1_122 gnd vdd FILL
XFILL_1_AOI21X1_11 gnd vdd FILL
XFILL_0_INVX1_133 gnd vdd FILL
XFILL_0_INVX1_144 gnd vdd FILL
XFILL_1_AOI21X1_22 gnd vdd FILL
XFILL_0_INVX1_155 gnd vdd FILL
XFILL_1_AOI21X1_33 gnd vdd FILL
XFILL_1_AOI21X1_44 gnd vdd FILL
XFILL_0_INVX1_166 gnd vdd FILL
XFILL_0_INVX1_177 gnd vdd FILL
XFILL_23_DFFSR_170 gnd vdd FILL
XFILL_1_AOI21X1_55 gnd vdd FILL
XFILL_11_OAI22X1_13 gnd vdd FILL
XFILL_60_6_0 gnd vdd FILL
XFILL_0_INVX1_188 gnd vdd FILL
XFILL_1_AOI21X1_66 gnd vdd FILL
XFILL_11_OAI22X1_24 gnd vdd FILL
XFILL_23_DFFSR_181 gnd vdd FILL
XFILL_0_INVX1_199 gnd vdd FILL
XFILL_4_INVX1_110 gnd vdd FILL
XFILL_1_AOI21X1_77 gnd vdd FILL
XFILL_32_3_2 gnd vdd FILL
XFILL_11_OAI22X1_35 gnd vdd FILL
XFILL_4_INVX1_121 gnd vdd FILL
XFILL_23_DFFSR_192 gnd vdd FILL
XFILL_11_OAI22X1_46 gnd vdd FILL
XFILL_4_INVX1_132 gnd vdd FILL
XFILL_4_NOR2X1_110 gnd vdd FILL
XFILL_15_OAI21X1_15 gnd vdd FILL
XFILL_4_INVX1_143 gnd vdd FILL
XFILL_4_NOR2X1_121 gnd vdd FILL
XFILL_15_OAI21X1_26 gnd vdd FILL
XFILL_4_INVX1_154 gnd vdd FILL
XFILL_4_NOR2X1_132 gnd vdd FILL
XFILL_4_INVX1_165 gnd vdd FILL
XFILL_15_OAI21X1_37 gnd vdd FILL
XFILL_4_NOR2X1_143 gnd vdd FILL
XFILL_15_OAI21X1_48 gnd vdd FILL
XFILL_4_INVX1_176 gnd vdd FILL
XFILL_4_NOR2X1_154 gnd vdd FILL
XFILL_27_DFFSR_180 gnd vdd FILL
XFILL_4_NOR2X1_165 gnd vdd FILL
XFILL_4_INVX1_187 gnd vdd FILL
XFILL_4_NOR2X1_176 gnd vdd FILL
XFILL_4_INVX1_198 gnd vdd FILL
XFILL_27_DFFSR_191 gnd vdd FILL
XFILL_4_NOR2X1_187 gnd vdd FILL
XFILL_4_NOR2X1_198 gnd vdd FILL
XFILL_21_MUX2X1_101 gnd vdd FILL
XFILL_21_MUX2X1_112 gnd vdd FILL
XFILL_21_MUX2X1_123 gnd vdd FILL
XFILL_2_OAI22X1_5 gnd vdd FILL
XFILL_21_MUX2X1_134 gnd vdd FILL
XFILL_21_MUX2X1_145 gnd vdd FILL
XFILL_21_MUX2X1_156 gnd vdd FILL
XFILL_60_15 gnd vdd FILL
XFILL_21_MUX2X1_167 gnd vdd FILL
XFILL_73_DFFSR_270 gnd vdd FILL
XFILL_21_MUX2X1_178 gnd vdd FILL
XFILL_4_MUX2X1_105 gnd vdd FILL
XFILL_21_MUX2X1_189 gnd vdd FILL
XFILL_4_MUX2X1_116 gnd vdd FILL
XFILL_4_MUX2X1_127 gnd vdd FILL
XFILL_4_MUX2X1_138 gnd vdd FILL
XFILL_4_MUX2X1_149 gnd vdd FILL
XFILL_6_OAI22X1_4 gnd vdd FILL
XFILL_1_OAI22X1_30 gnd vdd FILL
XFILL_1_OAI22X1_41 gnd vdd FILL
XFILL_5_OAI21X1_10 gnd vdd FILL
XFILL_5_OAI21X1_21 gnd vdd FILL
XFILL_5_OAI21X1_32 gnd vdd FILL
XFILL_51_DFFSR_205 gnd vdd FILL
XFILL_51_DFFSR_216 gnd vdd FILL
XFILL_5_OAI21X1_43 gnd vdd FILL
XFILL_51_DFFSR_227 gnd vdd FILL
XFILL_51_DFFSR_238 gnd vdd FILL
XFILL_51_DFFSR_249 gnd vdd FILL
XFILL_5_DFFSR_4 gnd vdd FILL
XFILL_55_DFFSR_204 gnd vdd FILL
XFILL_55_DFFSR_215 gnd vdd FILL
XFILL_51_6_0 gnd vdd FILL
XFILL_18_DFFSR_2 gnd vdd FILL
XFILL_55_DFFSR_226 gnd vdd FILL
XFILL_23_3_2 gnd vdd FILL
XFILL_75_DFFSR_3 gnd vdd FILL
XFILL_55_DFFSR_237 gnd vdd FILL
XFILL_9_BUFX4_12 gnd vdd FILL
XFILL_55_DFFSR_248 gnd vdd FILL
XFILL_11_NAND3X1_106 gnd vdd FILL
XFILL_9_BUFX4_23 gnd vdd FILL
XFILL_11_NAND3X1_117 gnd vdd FILL
XFILL_11_NAND3X1_128 gnd vdd FILL
XFILL_55_DFFSR_259 gnd vdd FILL
XFILL_9_BUFX4_34 gnd vdd FILL
XFILL_9_BUFX4_45 gnd vdd FILL
XFILL_82_DFFSR_104 gnd vdd FILL
XFILL_59_DFFSR_203 gnd vdd FILL
XFILL_9_BUFX4_56 gnd vdd FILL
XFILL_82_DFFSR_115 gnd vdd FILL
XFILL_9_BUFX4_67 gnd vdd FILL
XFILL_9_BUFX4_78 gnd vdd FILL
XFILL_82_DFFSR_126 gnd vdd FILL
XFILL_59_DFFSR_214 gnd vdd FILL
XFILL_59_DFFSR_225 gnd vdd FILL
XFILL_9_BUFX4_89 gnd vdd FILL
XFILL_82_DFFSR_137 gnd vdd FILL
XFILL_59_DFFSR_236 gnd vdd FILL
XFILL_82_DFFSR_148 gnd vdd FILL
XFILL_59_DFFSR_247 gnd vdd FILL
XFILL_59_DFFSR_258 gnd vdd FILL
XFILL_82_DFFSR_159 gnd vdd FILL
XFILL_59_DFFSR_269 gnd vdd FILL
XFILL_2_DFFSR_207 gnd vdd FILL
XFILL_86_DFFSR_103 gnd vdd FILL
XFILL_86_DFFSR_114 gnd vdd FILL
XFILL_2_DFFSR_218 gnd vdd FILL
XFILL_7_NAND3X1_19 gnd vdd FILL
XFILL_2_DFFSR_229 gnd vdd FILL
XFILL_86_DFFSR_125 gnd vdd FILL
XFILL_86_DFFSR_136 gnd vdd FILL
XFILL_86_DFFSR_147 gnd vdd FILL
XFILL_86_DFFSR_158 gnd vdd FILL
XFILL_10_BUFX4_105 gnd vdd FILL
XFILL_86_DFFSR_169 gnd vdd FILL
XFILL_18_CLKBUF1_9 gnd vdd FILL
XFILL_6_DFFSR_206 gnd vdd FILL
XFILL_3_NAND3X1_6 gnd vdd FILL
XFILL_6_DFFSR_217 gnd vdd FILL
XFILL_6_DFFSR_228 gnd vdd FILL
XFILL_10_NOR2X1_190 gnd vdd FILL
XFILL_6_DFFSR_239 gnd vdd FILL
XFILL_53_DFFSR_19 gnd vdd FILL
XFILL_14_BUFX4_104 gnd vdd FILL
XFILL_59_7_0 gnd vdd FILL
XFILL_40_DFFSR_270 gnd vdd FILL
XFILL_6_4_2 gnd vdd FILL
XFILL_7_NAND3X1_5 gnd vdd FILL
XMUX2X1_19 BUFX4_71/Y INVX1_32/Y MUX2X1_20/S gnd DFFSR_12/D vdd MUX2X1
XFILL_12_BUFX4_2 gnd vdd FILL
XFILL_22_DFFSR_18 gnd vdd FILL
XFILL_13_BUFX4_50 gnd vdd FILL
XFILL_22_DFFSR_29 gnd vdd FILL
XFILL_13_BUFX4_61 gnd vdd FILL
XFILL_13_BUFX4_72 gnd vdd FILL
XFILL_10_MUX2X1_130 gnd vdd FILL
XFILL_13_BUFX4_83 gnd vdd FILL
XFILL_10_MUX2X1_141 gnd vdd FILL
XFILL_10_MUX2X1_152 gnd vdd FILL
XFILL_13_BUFX4_94 gnd vdd FILL
XFILL_10_MUX2X1_163 gnd vdd FILL
XFILL_71_DFFSR_180 gnd vdd FILL
XFILL_42_6_0 gnd vdd FILL
XFILL_10_MUX2X1_174 gnd vdd FILL
XFILL_10_MUX2X1_185 gnd vdd FILL
XFILL_14_3_2 gnd vdd FILL
XFILL_62_DFFSR_17 gnd vdd FILL
XFILL_71_DFFSR_191 gnd vdd FILL
XFILL_62_DFFSR_28 gnd vdd FILL
XFILL_22_DFFSR_204 gnd vdd FILL
XFILL_22_DFFSR_215 gnd vdd FILL
XFILL_62_DFFSR_39 gnd vdd FILL
XFILL_22_DFFSR_226 gnd vdd FILL
XFILL_22_DFFSR_237 gnd vdd FILL
XFILL_22_DFFSR_248 gnd vdd FILL
XFILL_22_DFFSR_259 gnd vdd FILL
XFILL_75_DFFSR_190 gnd vdd FILL
XFILL_26_DFFSR_203 gnd vdd FILL
XAOI22X1_2 OAI21X1_1/C AOI22X1_3/A AOI22X1_2/C AOI22X1_2/D gnd AND2X2_2/B vdd AOI22X1
XFILL_5_DFFSR_19 gnd vdd FILL
XFILL_26_DFFSR_214 gnd vdd FILL
XFILL_26_DFFSR_225 gnd vdd FILL
XFILL_31_DFFSR_16 gnd vdd FILL
XFILL_26_DFFSR_236 gnd vdd FILL
XFILL_26_DFFSR_247 gnd vdd FILL
XFILL_31_DFFSR_27 gnd vdd FILL
XFILL_31_DFFSR_38 gnd vdd FILL
XFILL_26_DFFSR_258 gnd vdd FILL
XINVX1_201 DFFSR_85/Q gnd INVX1_201/Y vdd INVX1
XFILL_26_DFFSR_269 gnd vdd FILL
XINVX1_212 DFFSR_73/Q gnd INVX1_212/Y vdd INVX1
XFILL_31_DFFSR_49 gnd vdd FILL
XFILL_7_INVX1_40 gnd vdd FILL
XFILL_7_INVX1_51 gnd vdd FILL
XFILL_7_INVX1_209 gnd vdd FILL
XFILL_53_DFFSR_103 gnd vdd FILL
XINVX1_223 DFFSR_66/Q gnd INVX1_223/Y vdd INVX1
XFILL_7_INVX1_62 gnd vdd FILL
XFILL_53_DFFSR_114 gnd vdd FILL
XFILL_7_INVX1_73 gnd vdd FILL
XFILL_53_DFFSR_125 gnd vdd FILL
XFILL_7_INVX1_84 gnd vdd FILL
XFILL_53_DFFSR_136 gnd vdd FILL
XFILL_7_INVX1_95 gnd vdd FILL
XFILL_71_DFFSR_15 gnd vdd FILL
XFILL_71_DFFSR_26 gnd vdd FILL
XFILL_53_DFFSR_147 gnd vdd FILL
XFILL_53_DFFSR_158 gnd vdd FILL
XFILL_71_DFFSR_37 gnd vdd FILL
XFILL_53_DFFSR_169 gnd vdd FILL
XFILL_14_MUX2X1_5 gnd vdd FILL
XFILL_71_DFFSR_48 gnd vdd FILL
XFILL_71_DFFSR_59 gnd vdd FILL
XFILL_57_DFFSR_102 gnd vdd FILL
XFILL_57_DFFSR_113 gnd vdd FILL
XFILL_57_DFFSR_124 gnd vdd FILL
XFILL_7_NOR2X1_109 gnd vdd FILL
XFILL_57_DFFSR_135 gnd vdd FILL
XFILL_57_DFFSR_146 gnd vdd FILL
XFILL_13_NAND3X1_11 gnd vdd FILL
XNAND2X1_12 INVX1_218/A NOR2X1_13/Y gnd NOR2X1_68/A vdd NAND2X1
XFILL_57_DFFSR_157 gnd vdd FILL
XFILL_13_NAND3X1_22 gnd vdd FILL
XNAND2X1_23 INVX4_1/A INVX1_205/A gnd NAND2X1_23/Y vdd NAND2X1
XFILL_57_DFFSR_168 gnd vdd FILL
XFILL_13_NAND3X1_33 gnd vdd FILL
XFILL_0_MUX2X1_180 gnd vdd FILL
XNAND2X1_34 INVX1_141/Y NOR2X1_122/Y gnd OR2X2_1/B vdd NAND2X1
XFILL_57_DFFSR_179 gnd vdd FILL
XFILL_2_INVX8_2 gnd vdd FILL
XFILL_13_NAND3X1_44 gnd vdd FILL
XNAND2X1_45 NOR2X1_1/Y NOR2X1_122/Y gnd NOR2X1_25/A vdd NAND2X1
XFILL_0_MUX2X1_191 gnd vdd FILL
XFILL_0_DFFSR_106 gnd vdd FILL
XFILL_13_NAND3X1_55 gnd vdd FILL
XFILL_5_BUFX4_60 gnd vdd FILL
XFILL_40_DFFSR_14 gnd vdd FILL
XFILL_5_BUFX4_71 gnd vdd FILL
XFILL_0_DFFSR_117 gnd vdd FILL
XFILL_40_DFFSR_25 gnd vdd FILL
XNAND2X1_56 INVX1_218/A NOR2X1_122/Y gnd NOR2X1_27/A vdd NAND2X1
XFILL_33_CLKBUF1_11 gnd vdd FILL
XFILL_13_NAND3X1_66 gnd vdd FILL
XFILL_40_DFFSR_36 gnd vdd FILL
XFILL_5_BUFX4_82 gnd vdd FILL
XNAND2X1_67 INVX1_57/A NOR2X1_122/Y gnd NOR2X1_7/A vdd NAND2X1
XFILL_33_CLKBUF1_22 gnd vdd FILL
XFILL_13_NAND3X1_77 gnd vdd FILL
XNAND2X1_78 INVX4_1/A INVX1_160/Y gnd NAND2X1_78/Y vdd NAND2X1
XFILL_5_BUFX4_93 gnd vdd FILL
XFILL_0_DFFSR_128 gnd vdd FILL
XFILL_13_NAND3X1_88 gnd vdd FILL
XFILL_33_CLKBUF1_33 gnd vdd FILL
XNAND2X1_89 INVX4_1/A INVX1_3/A gnd NAND2X1_89/Y vdd NAND2X1
XFILL_0_DFFSR_139 gnd vdd FILL
XFILL_40_DFFSR_47 gnd vdd FILL
XFILL_13_NAND3X1_99 gnd vdd FILL
XFILL_40_DFFSR_58 gnd vdd FILL
XFILL_64_2_2 gnd vdd FILL
XFILL_40_DFFSR_69 gnd vdd FILL
XFILL_42_4 gnd vdd FILL
XFILL_80_DFFSR_13 gnd vdd FILL
XFILL_4_DFFSR_105 gnd vdd FILL
XFILL_80_DFFSR_24 gnd vdd FILL
XFILL_4_DFFSR_116 gnd vdd FILL
XFILL_80_DFFSR_35 gnd vdd FILL
XFILL_4_DFFSR_127 gnd vdd FILL
XFILL_80_DFFSR_46 gnd vdd FILL
XFILL_4_DFFSR_138 gnd vdd FILL
XFILL_23_MUX2X1_3 gnd vdd FILL
XFILL_4_DFFSR_149 gnd vdd FILL
XFILL_80_DFFSR_57 gnd vdd FILL
XFILL_33_6_0 gnd vdd FILL
XFILL_80_DFFSR_68 gnd vdd FILL
XFILL_80_DFFSR_79 gnd vdd FILL
XFILL_28_2 gnd vdd FILL
XFILL_8_DFFSR_104 gnd vdd FILL
XFILL_7_NOR2X1_6 gnd vdd FILL
XFILL_12_MUX2X1_13 gnd vdd FILL
XFILL_8_DFFSR_115 gnd vdd FILL
XFILL_8_DFFSR_126 gnd vdd FILL
XFILL_12_MUX2X1_24 gnd vdd FILL
XFILL_8_DFFSR_137 gnd vdd FILL
XFILL_12_MUX2X1_35 gnd vdd FILL
XFILL_8_DFFSR_148 gnd vdd FILL
XFILL_12_MUX2X1_46 gnd vdd FILL
XFILL_8_DFFSR_159 gnd vdd FILL
XFILL_12_MUX2X1_57 gnd vdd FILL
XAOI22X1_10 AND2X2_4/Y NOR2X1_6/A DFFSR_5/Q INVX1_123/Y gnd NAND3X1_17/A vdd AOI22X1
XFILL_4_OAI22X1_18 gnd vdd FILL
XFILL_12_MUX2X1_68 gnd vdd FILL
XFILL_12_MUX2X1_79 gnd vdd FILL
XFILL_20_NOR3X1_9 gnd vdd FILL
XFILL_4_OAI22X1_29 gnd vdd FILL
XFILL_0_NOR3X1_17 gnd vdd FILL
XFILL_0_NOR3X1_28 gnd vdd FILL
XFILL_42_DFFSR_190 gnd vdd FILL
XFILL_0_NOR3X1_39 gnd vdd FILL
XFILL_16_MUX2X1_12 gnd vdd FILL
XFILL_16_MUX2X1_23 gnd vdd FILL
XFILL_17_AOI22X1_11 gnd vdd FILL
XFILL_16_MUX2X1_34 gnd vdd FILL
XFILL_16_MUX2X1_45 gnd vdd FILL
XFILL_6_MUX2X1_4 gnd vdd FILL
XFILL_16_MUX2X1_56 gnd vdd FILL
XFILL_16_MUX2X1_67 gnd vdd FILL
XFILL_16_MUX2X1_78 gnd vdd FILL
XFILL_3_NAND3X1_50 gnd vdd FILL
XFILL_4_NOR3X1_16 gnd vdd FILL
XFILL_3_NAND3X1_61 gnd vdd FILL
XFILL_16_MUX2X1_89 gnd vdd FILL
XFILL_4_NOR3X1_27 gnd vdd FILL
XFILL_3_NAND3X1_72 gnd vdd FILL
XFILL_41_DFFSR_6 gnd vdd FILL
XFILL_4_NOR3X1_38 gnd vdd FILL
XFILL_7_NAND2X1_30 gnd vdd FILL
XFILL_9_DFFSR_5 gnd vdd FILL
XFILL_4_NOR3X1_49 gnd vdd FILL
XFILL_20_DFFSR_103 gnd vdd FILL
XFILL_7_NAND2X1_41 gnd vdd FILL
XFILL_3_NAND3X1_83 gnd vdd FILL
XFILL_3_NAND3X1_94 gnd vdd FILL
XFILL_7_NAND2X1_52 gnd vdd FILL
XFILL_20_DFFSR_114 gnd vdd FILL
XFILL_20_DFFSR_125 gnd vdd FILL
XFILL_7_NAND2X1_63 gnd vdd FILL
XFILL_20_DFFSR_136 gnd vdd FILL
XFILL_79_DFFSR_4 gnd vdd FILL
XFILL_7_NAND2X1_74 gnd vdd FILL
XFILL_7_NAND2X1_85 gnd vdd FILL
XFILL_20_DFFSR_147 gnd vdd FILL
XFILL_20_DFFSR_158 gnd vdd FILL
XFILL_8_NOR3X1_15 gnd vdd FILL
XFILL_7_NAND2X1_96 gnd vdd FILL
XFILL_20_DFFSR_169 gnd vdd FILL
XFILL_8_NOR3X1_26 gnd vdd FILL
XFILL_1_INVX1_109 gnd vdd FILL
XFILL_8_NOR3X1_37 gnd vdd FILL
XFILL_24_DFFSR_102 gnd vdd FILL
XFILL_8_NOR3X1_48 gnd vdd FILL
XFILL_15_CLKBUF1_16 gnd vdd FILL
XFILL_24_DFFSR_113 gnd vdd FILL
XFILL_24_DFFSR_124 gnd vdd FILL
XFILL_15_CLKBUF1_27 gnd vdd FILL
XFILL_15_CLKBUF1_38 gnd vdd FILL
XFILL_24_DFFSR_135 gnd vdd FILL
XFILL_24_DFFSR_146 gnd vdd FILL
XFILL_10_AOI21X1_13 gnd vdd FILL
XFILL_24_DFFSR_157 gnd vdd FILL
XFILL_10_AOI21X1_24 gnd vdd FILL
XFILL_24_DFFSR_168 gnd vdd FILL
XFILL_10_AOI21X1_35 gnd vdd FILL
XFILL_24_DFFSR_179 gnd vdd FILL
XFILL_10_AOI21X1_46 gnd vdd FILL
XFILL_5_INVX1_108 gnd vdd FILL
XFILL_1_DFFSR_12 gnd vdd FILL
XFILL_55_2_2 gnd vdd FILL
XFILL_28_DFFSR_101 gnd vdd FILL
XFILL_10_AOI21X1_57 gnd vdd FILL
XFILL_5_INVX1_119 gnd vdd FILL
XFILL_10_AOI21X1_68 gnd vdd FILL
XFILL_1_DFFSR_23 gnd vdd FILL
XFILL_28_DFFSR_112 gnd vdd FILL
XFILL_1_DFFSR_34 gnd vdd FILL
XFILL_10_AOI21X1_79 gnd vdd FILL
XFILL_28_DFFSR_123 gnd vdd FILL
XFILL_28_DFFSR_134 gnd vdd FILL
XFILL_1_DFFSR_45 gnd vdd FILL
XFILL_1_DFFSR_56 gnd vdd FILL
XFILL_28_DFFSR_145 gnd vdd FILL
XFILL_1_DFFSR_67 gnd vdd FILL
XFILL_28_DFFSR_156 gnd vdd FILL
XFILL_1_DFFSR_78 gnd vdd FILL
XFILL_28_DFFSR_167 gnd vdd FILL
XFILL_1_DFFSR_89 gnd vdd FILL
XFILL_28_DFFSR_178 gnd vdd FILL
XFILL_20_NOR3X1_14 gnd vdd FILL
XFILL_28_DFFSR_189 gnd vdd FILL
XFILL_24_6_0 gnd vdd FILL
XFILL_20_NOR3X1_25 gnd vdd FILL
XFILL_20_NOR3X1_36 gnd vdd FILL
XFILL_20_NOR3X1_47 gnd vdd FILL
XFILL_70_DFFSR_203 gnd vdd FILL
XFILL_70_DFFSR_214 gnd vdd FILL
XFILL_70_DFFSR_225 gnd vdd FILL
XFILL_70_DFFSR_236 gnd vdd FILL
XFILL_12_NAND3X1_107 gnd vdd FILL
XFILL_70_DFFSR_247 gnd vdd FILL
XFILL_49_DFFSR_80 gnd vdd FILL
XFILL_24_NOR3X1_13 gnd vdd FILL
XFILL_12_NAND3X1_118 gnd vdd FILL
XFILL_12_NAND3X1_129 gnd vdd FILL
XFILL_49_DFFSR_91 gnd vdd FILL
XFILL_70_DFFSR_258 gnd vdd FILL
XFILL_70_DFFSR_269 gnd vdd FILL
XFILL_24_NOR3X1_24 gnd vdd FILL
XFILL_24_NOR3X1_35 gnd vdd FILL
XFILL_74_DFFSR_202 gnd vdd FILL
XFILL_24_NOR3X1_46 gnd vdd FILL
XFILL_74_DFFSR_213 gnd vdd FILL
XFILL_22_CLKBUF1_40 gnd vdd FILL
XFILL_74_DFFSR_224 gnd vdd FILL
XFILL_74_DFFSR_235 gnd vdd FILL
XFILL_74_DFFSR_246 gnd vdd FILL
XFILL_5_CLKBUF1_11 gnd vdd FILL
XFILL_28_NOR3X1_12 gnd vdd FILL
XFILL_74_DFFSR_257 gnd vdd FILL
XFILL_3_BUFX4_5 gnd vdd FILL
XFILL_28_NOR3X1_23 gnd vdd FILL
XFILL_5_CLKBUF1_22 gnd vdd FILL
XFILL_74_DFFSR_268 gnd vdd FILL
XFILL_28_NOR3X1_34 gnd vdd FILL
XFILL_5_CLKBUF1_33 gnd vdd FILL
XFILL_78_DFFSR_201 gnd vdd FILL
XFILL_28_NOR3X1_45 gnd vdd FILL
XOAI22X1_5 OAI22X1_5/A OAI22X1_5/B INVX1_7/Y OAI22X1_5/D gnd OAI22X1_5/Y vdd OAI22X1
XFILL_78_DFFSR_212 gnd vdd FILL
XFILL_13_MUX2X1_107 gnd vdd FILL
XFILL_18_DFFSR_90 gnd vdd FILL
XFILL_13_MUX2X1_118 gnd vdd FILL
XFILL_13_MUX2X1_129 gnd vdd FILL
XFILL_0_AOI21X1_30 gnd vdd FILL
XFILL_78_DFFSR_223 gnd vdd FILL
XFILL_78_DFFSR_234 gnd vdd FILL
XFILL_0_AOI21X1_41 gnd vdd FILL
XFILL_0_AOI21X1_52 gnd vdd FILL
XFILL_78_DFFSR_245 gnd vdd FILL
XFILL_78_DFFSR_256 gnd vdd FILL
XFILL_10_OAI22X1_10 gnd vdd FILL
XFILL_0_AOI21X1_63 gnd vdd FILL
XFILL_10_OAI22X1_21 gnd vdd FILL
XFILL_0_AOI21X1_74 gnd vdd FILL
XFILL_78_DFFSR_267 gnd vdd FILL
XFILL_33_CLKBUF1_8 gnd vdd FILL
XFILL_10_OAI22X1_32 gnd vdd FILL
XFILL_10_OAI22X1_43 gnd vdd FILL
XFILL_14_OAI21X1_12 gnd vdd FILL
XFILL_14_OAI21X1_23 gnd vdd FILL
XFILL_7_7_0 gnd vdd FILL
XFILL_3_NOR2X1_140 gnd vdd FILL
XFILL_14_OAI21X1_34 gnd vdd FILL
XFILL_14_OAI21X1_45 gnd vdd FILL
XFILL_3_NOR2X1_151 gnd vdd FILL
XFILL_3_NOR2X1_162 gnd vdd FILL
XFILL_3_NOR2X1_173 gnd vdd FILL
XFILL_2_INVX1_9 gnd vdd FILL
XFILL_3_NOR2X1_184 gnd vdd FILL
XFILL_3_NOR2X1_195 gnd vdd FILL
XFILL_46_2_2 gnd vdd FILL
XFILL_20_MUX2X1_120 gnd vdd FILL
XFILL_15_6_0 gnd vdd FILL
XFILL_20_MUX2X1_131 gnd vdd FILL
XFILL_20_MUX2X1_142 gnd vdd FILL
XFILL_20_MUX2X1_153 gnd vdd FILL
XFILL_21_9 gnd vdd FILL
XFILL_3_MUX2X1_102 gnd vdd FILL
XFILL_20_MUX2X1_164 gnd vdd FILL
XFILL_20_MUX2X1_175 gnd vdd FILL
XFILL_3_MUX2X1_113 gnd vdd FILL
XFILL_20_MUX2X1_186 gnd vdd FILL
XFILL_3_MUX2X1_124 gnd vdd FILL
XFILL_14_8 gnd vdd FILL
XFILL_3_MUX2X1_135 gnd vdd FILL
XFILL_3_MUX2X1_146 gnd vdd FILL
XFILL_14_BUFX4_17 gnd vdd FILL
XFILL_3_MUX2X1_157 gnd vdd FILL
XFILL_14_BUFX4_28 gnd vdd FILL
XFILL_3_MUX2X1_168 gnd vdd FILL
XFILL_14_BUFX4_39 gnd vdd FILL
XFILL_3_MUX2X1_179 gnd vdd FILL
XFILL_6_INVX8_3 gnd vdd FILL
XDFFSR_207 NOR2X1_26/A CLKBUF1_4/Y DFFSR_90/R vdd DFFSR_207/D gnd vdd DFFSR
XDFFSR_218 INVX1_76/A DFFSR_7/CLK DFFSR_26/R vdd MUX2X1_63/Y gnd vdd DFFSR
XFILL_19_INVX8_1 gnd vdd FILL
XDFFSR_229 INVX1_70/A DFFSR_7/CLK DFFSR_26/R vdd MUX2X1_56/Y gnd vdd DFFSR
XFILL_41_DFFSR_202 gnd vdd FILL
XFILL_4_OAI21X1_40 gnd vdd FILL
XFILL_41_DFFSR_213 gnd vdd FILL
XFILL_3_OAI21X1_3 gnd vdd FILL
XFILL_41_DFFSR_224 gnd vdd FILL
XFILL_41_DFFSR_235 gnd vdd FILL
XFILL_41_DFFSR_246 gnd vdd FILL
XFILL_0_NOR2X1_50 gnd vdd FILL
XFILL_0_NOR2X1_61 gnd vdd FILL
XFILL_41_DFFSR_257 gnd vdd FILL
XFILL_0_NOR2X1_72 gnd vdd FILL
XFILL_41_DFFSR_268 gnd vdd FILL
XFILL_0_NOR2X1_83 gnd vdd FILL
XFILL_0_NOR2X1_94 gnd vdd FILL
XFILL_45_DFFSR_201 gnd vdd FILL
XFILL_23_DFFSR_3 gnd vdd FILL
XFILL_7_OAI21X1_2 gnd vdd FILL
XFILL_45_DFFSR_212 gnd vdd FILL
XFILL_80_DFFSR_4 gnd vdd FILL
XFILL_45_DFFSR_223 gnd vdd FILL
XFILL_45_DFFSR_234 gnd vdd FILL
XFILL_45_DFFSR_245 gnd vdd FILL
XFILL_4_NOR2X1_60 gnd vdd FILL
XFILL_45_DFFSR_256 gnd vdd FILL
XFILL_4_NOR2X1_71 gnd vdd FILL
XFILL_45_DFFSR_267 gnd vdd FILL
XFILL_4_NOR2X1_82 gnd vdd FILL
XFILL_4_NOR2X1_93 gnd vdd FILL
XFILL_72_DFFSR_101 gnd vdd FILL
XFILL_49_DFFSR_200 gnd vdd FILL
XFILL_49_DFFSR_211 gnd vdd FILL
XFILL_72_DFFSR_112 gnd vdd FILL
XFILL_72_DFFSR_123 gnd vdd FILL
XFILL_72_DFFSR_134 gnd vdd FILL
XFILL_49_DFFSR_222 gnd vdd FILL
XFILL_49_DFFSR_233 gnd vdd FILL
XFILL_72_DFFSR_145 gnd vdd FILL
XFILL_49_DFFSR_244 gnd vdd FILL
XFILL_72_DFFSR_156 gnd vdd FILL
XFILL_49_DFFSR_255 gnd vdd FILL
XFILL_72_DFFSR_167 gnd vdd FILL
XFILL_8_NOR2X1_70 gnd vdd FILL
XFILL_49_DFFSR_266 gnd vdd FILL
XFILL_72_DFFSR_178 gnd vdd FILL
XFILL_8_NOR2X1_81 gnd vdd FILL
XFILL_65_5_0 gnd vdd FILL
XFILL_8_NOR2X1_92 gnd vdd FILL
XFILL_72_DFFSR_189 gnd vdd FILL
XFILL_76_DFFSR_100 gnd vdd FILL
XFILL_37_2_2 gnd vdd FILL
XFILL_76_DFFSR_111 gnd vdd FILL
XFILL_6_NAND3X1_16 gnd vdd FILL
XFILL_76_DFFSR_122 gnd vdd FILL
XFILL_76_DFFSR_133 gnd vdd FILL
XFILL_6_NAND3X1_27 gnd vdd FILL
XFILL_76_DFFSR_144 gnd vdd FILL
XFILL_6_NAND3X1_38 gnd vdd FILL
XFILL_76_DFFSR_155 gnd vdd FILL
XFILL_6_NAND3X1_49 gnd vdd FILL
XFILL_76_DFFSR_166 gnd vdd FILL
XFILL_76_DFFSR_177 gnd vdd FILL
XFILL_45_DFFSR_7 gnd vdd FILL
XFILL_6_BUFX4_16 gnd vdd FILL
XFILL_76_DFFSR_188 gnd vdd FILL
XFILL_6_BUFX4_27 gnd vdd FILL
XFILL_76_DFFSR_199 gnd vdd FILL
XFILL_6_BUFX4_38 gnd vdd FILL
XFILL_6_BUFX4_49 gnd vdd FILL
XFILL_0_NAND2X1_5 gnd vdd FILL
XFILL_20_1_2 gnd vdd FILL
XFILL_4_NAND2X1_4 gnd vdd FILL
XFILL_0_MUX2X1_90 gnd vdd FILL
XFILL_13_AND2X2_4 gnd vdd FILL
XFILL_8_NAND2X1_3 gnd vdd FILL
XFILL_12_DFFSR_201 gnd vdd FILL
XFILL_12_DFFSR_212 gnd vdd FILL
XFILL_12_DFFSR_223 gnd vdd FILL
XFILL_12_DFFSR_234 gnd vdd FILL
XFILL_12_DFFSR_245 gnd vdd FILL
XFILL_12_DFFSR_256 gnd vdd FILL
XFILL_12_DFFSR_267 gnd vdd FILL
XFILL_10_BUFX4_10 gnd vdd FILL
XFILL_16_DFFSR_200 gnd vdd FILL
XFILL_16_DFFSR_211 gnd vdd FILL
XFILL_10_BUFX4_21 gnd vdd FILL
XFILL_25_CLKBUF1_17 gnd vdd FILL
XFILL_25_CLKBUF1_28 gnd vdd FILL
XFILL_10_BUFX4_32 gnd vdd FILL
XFILL_16_DFFSR_222 gnd vdd FILL
XFILL_25_CLKBUF1_39 gnd vdd FILL
XFILL_56_5_0 gnd vdd FILL
XFILL_16_DFFSR_233 gnd vdd FILL
XFILL_10_BUFX4_43 gnd vdd FILL
XFILL_10_BUFX4_54 gnd vdd FILL
XFILL_16_DFFSR_244 gnd vdd FILL
XFILL_28_2_2 gnd vdd FILL
XFILL_16_DFFSR_255 gnd vdd FILL
XFILL_10_BUFX4_65 gnd vdd FILL
XFILL_3_2_2 gnd vdd FILL
XFILL_10_BUFX4_76 gnd vdd FILL
XFILL_7_BUFX4_6 gnd vdd FILL
XFILL_10_BUFX4_87 gnd vdd FILL
XFILL_16_DFFSR_266 gnd vdd FILL
XFILL_43_DFFSR_100 gnd vdd FILL
XFILL_10_BUFX4_98 gnd vdd FILL
XFILL_43_DFFSR_111 gnd vdd FILL
XFILL_43_DFFSR_122 gnd vdd FILL
XFILL_3_AOI21X1_18 gnd vdd FILL
XFILL_43_DFFSR_133 gnd vdd FILL
XFILL_4_AOI21X1_9 gnd vdd FILL
XFILL_3_AOI21X1_29 gnd vdd FILL
XFILL_43_DFFSR_144 gnd vdd FILL
XFILL_43_DFFSR_155 gnd vdd FILL
XFILL_43_DFFSR_166 gnd vdd FILL
XFILL_43_DFFSR_177 gnd vdd FILL
XFILL_43_DFFSR_188 gnd vdd FILL
XFILL_47_DFFSR_110 gnd vdd FILL
XFILL_43_DFFSR_199 gnd vdd FILL
XFILL_6_NOR2X1_106 gnd vdd FILL
XFILL_47_DFFSR_121 gnd vdd FILL
XFILL_47_DFFSR_132 gnd vdd FILL
XFILL_8_AOI21X1_8 gnd vdd FILL
XFILL_6_NOR2X1_117 gnd vdd FILL
XFILL_47_DFFSR_143 gnd vdd FILL
XFILL_6_NOR2X1_128 gnd vdd FILL
XFILL_6_NOR2X1_139 gnd vdd FILL
XFILL_47_DFFSR_154 gnd vdd FILL
XFILL_11_1_2 gnd vdd FILL
XFILL_13_NAND3X1_108 gnd vdd FILL
XFILL_47_DFFSR_165 gnd vdd FILL
XFILL_12_NAND3X1_30 gnd vdd FILL
XFILL_13_NAND3X1_119 gnd vdd FILL
XFILL_12_NAND3X1_41 gnd vdd FILL
XFILL_47_DFFSR_176 gnd vdd FILL
XFILL_4_INVX1_11 gnd vdd FILL
XFILL_47_DFFSR_187 gnd vdd FILL
XFILL_12_NAND3X1_52 gnd vdd FILL
XFILL_47_DFFSR_198 gnd vdd FILL
XFILL_4_INVX1_22 gnd vdd FILL
XFILL_12_NAND3X1_63 gnd vdd FILL
XFILL_4_INVX1_33 gnd vdd FILL
XFILL_12_NAND3X1_74 gnd vdd FILL
XFILL_4_INVX1_44 gnd vdd FILL
XFILL_5_AND2X2_3 gnd vdd FILL
XFILL_32_CLKBUF1_30 gnd vdd FILL
XFILL_12_NAND3X1_85 gnd vdd FILL
XFILL_4_INVX1_55 gnd vdd FILL
XFILL_32_CLKBUF1_41 gnd vdd FILL
XFILL_4_INVX1_66 gnd vdd FILL
XFILL_12_NAND3X1_96 gnd vdd FILL
XFILL_3_BUFX2_2 gnd vdd FILL
XFILL_4_INVX1_77 gnd vdd FILL
XFILL_13_AOI22X1_5 gnd vdd FILL
XFILL_4_INVX1_88 gnd vdd FILL
XFILL_4_INVX1_99 gnd vdd FILL
XFILL_11_MUX2X1_9 gnd vdd FILL
XFILL_23_MUX2X1_108 gnd vdd FILL
XFILL_23_MUX2X1_119 gnd vdd FILL
XFILL_17_AOI22X1_4 gnd vdd FILL
XFILL_2_BUFX4_20 gnd vdd FILL
XFILL_62_DFFSR_1 gnd vdd FILL
XFILL_2_BUFX4_31 gnd vdd FILL
XFILL_2_BUFX4_42 gnd vdd FILL
XFILL_19_DFFSR_13 gnd vdd FILL
XFILL_2_BUFX4_53 gnd vdd FILL
XFILL_19_DFFSR_24 gnd vdd FILL
XFILL_2_BUFX4_64 gnd vdd FILL
XFILL_19_DFFSR_35 gnd vdd FILL
XFILL_19_DFFSR_46 gnd vdd FILL
XFILL_2_BUFX4_75 gnd vdd FILL
XFILL_2_BUFX4_86 gnd vdd FILL
XFILL_2_BUFX4_97 gnd vdd FILL
XFILL_19_DFFSR_57 gnd vdd FILL
XFILL_3_OAI22X1_15 gnd vdd FILL
XFILL_19_DFFSR_68 gnd vdd FILL
XFILL_3_OAI22X1_26 gnd vdd FILL
XFILL_19_DFFSR_79 gnd vdd FILL
XFILL_3_OAI22X1_37 gnd vdd FILL
XFILL_3_OAI22X1_48 gnd vdd FILL
XFILL_47_5_0 gnd vdd FILL
XFILL_7_OAI21X1_17 gnd vdd FILL
XFILL_59_DFFSR_12 gnd vdd FILL
XFILL_7_OAI21X1_28 gnd vdd FILL
XFILL_19_2_2 gnd vdd FILL
XFILL_59_DFFSR_23 gnd vdd FILL
XFILL_59_DFFSR_34 gnd vdd FILL
XFILL_7_OAI21X1_39 gnd vdd FILL
XFILL_59_DFFSR_45 gnd vdd FILL
XFILL_59_DFFSR_56 gnd vdd FILL
XFILL_59_DFFSR_67 gnd vdd FILL
XFILL_20_MUX2X1_7 gnd vdd FILL
XFILL_59_DFFSR_78 gnd vdd FILL
XFILL_59_DFFSR_89 gnd vdd FILL
XFILL_2_NAND3X1_80 gnd vdd FILL
XFILL_10_DFFSR_100 gnd vdd FILL
XFILL_27_DFFSR_4 gnd vdd FILL
XFILL_61_0_2 gnd vdd FILL
XFILL_2_NAND3X1_91 gnd vdd FILL
XFILL_10_DFFSR_111 gnd vdd FILL
XFILL_6_NAND2X1_60 gnd vdd FILL
XFILL_0_NOR2X1_206 gnd vdd FILL
XFILL_10_DFFSR_122 gnd vdd FILL
XFILL_10_DFFSR_133 gnd vdd FILL
XFILL_84_DFFSR_5 gnd vdd FILL
XFILL_28_DFFSR_11 gnd vdd FILL
XFILL_6_NAND2X1_71 gnd vdd FILL
XFILL_10_DFFSR_144 gnd vdd FILL
XFILL_6_NAND2X1_82 gnd vdd FILL
XFILL_10_DFFSR_155 gnd vdd FILL
XFILL_28_DFFSR_22 gnd vdd FILL
XFILL_6_NAND2X1_93 gnd vdd FILL
XFILL_10_DFFSR_166 gnd vdd FILL
XFILL_28_DFFSR_33 gnd vdd FILL
XFILL_10_DFFSR_177 gnd vdd FILL
XFILL_3_INVX2_2 gnd vdd FILL
XFILL_28_DFFSR_44 gnd vdd FILL
XFILL_28_DFFSR_55 gnd vdd FILL
XFILL_12_5 gnd vdd FILL
XFILL_28_DFFSR_66 gnd vdd FILL
XFILL_10_DFFSR_188 gnd vdd FILL
XFILL_30_4_0 gnd vdd FILL
XFILL_14_DFFSR_110 gnd vdd FILL
XFILL_10_DFFSR_199 gnd vdd FILL
XFILL_14_CLKBUF1_13 gnd vdd FILL
XFILL_28_DFFSR_77 gnd vdd FILL
XFILL_14_CLKBUF1_24 gnd vdd FILL
XFILL_14_DFFSR_121 gnd vdd FILL
XFILL_14_DFFSR_132 gnd vdd FILL
XFILL_14_CLKBUF1_35 gnd vdd FILL
XFILL_28_DFFSR_88 gnd vdd FILL
XFILL_14_DFFSR_143 gnd vdd FILL
XFILL_28_DFFSR_99 gnd vdd FILL
XFILL_68_DFFSR_10 gnd vdd FILL
XFILL_68_DFFSR_21 gnd vdd FILL
XFILL_14_DFFSR_154 gnd vdd FILL
XFILL_14_DFFSR_165 gnd vdd FILL
XFILL_68_DFFSR_32 gnd vdd FILL
XFILL_68_DFFSR_43 gnd vdd FILL
XFILL_3_MUX2X1_8 gnd vdd FILL
XFILL_3_CLKBUF1_8 gnd vdd FILL
XFILL_14_DFFSR_176 gnd vdd FILL
XFILL_14_DFFSR_187 gnd vdd FILL
XFILL_68_DFFSR_54 gnd vdd FILL
XFILL_68_DFFSR_65 gnd vdd FILL
XFILL_68_DFFSR_76 gnd vdd FILL
XFILL_14_DFFSR_198 gnd vdd FILL
XFILL_18_DFFSR_120 gnd vdd FILL
XFILL_18_DFFSR_131 gnd vdd FILL
XFILL_68_DFFSR_87 gnd vdd FILL
XFILL_68_DFFSR_98 gnd vdd FILL
XFILL_18_DFFSR_142 gnd vdd FILL
XFILL_18_DFFSR_153 gnd vdd FILL
XFILL_18_DFFSR_164 gnd vdd FILL
XFILL_7_CLKBUF1_7 gnd vdd FILL
XFILL_10_NOR3X1_11 gnd vdd FILL
XFILL_18_DFFSR_175 gnd vdd FILL
XFILL_49_DFFSR_8 gnd vdd FILL
XFILL_18_DFFSR_186 gnd vdd FILL
XFILL_18_DFFSR_197 gnd vdd FILL
XFILL_37_DFFSR_20 gnd vdd FILL
XFILL_10_NOR3X1_22 gnd vdd FILL
XFILL_10_NOR3X1_33 gnd vdd FILL
XFILL_37_DFFSR_31 gnd vdd FILL
XFILL_60_DFFSR_200 gnd vdd FILL
XFILL_10_NOR3X1_44 gnd vdd FILL
XFILL_37_DFFSR_42 gnd vdd FILL
XFILL_60_DFFSR_211 gnd vdd FILL
XFILL_37_DFFSR_53 gnd vdd FILL
XFILL_60_DFFSR_222 gnd vdd FILL
XFILL_37_DFFSR_64 gnd vdd FILL
XFILL_60_DFFSR_233 gnd vdd FILL
XFILL_3_BUFX4_102 gnd vdd FILL
XFILL_37_DFFSR_75 gnd vdd FILL
XFILL_37_DFFSR_86 gnd vdd FILL
XFILL_60_DFFSR_244 gnd vdd FILL
XFILL_14_NOR3X1_10 gnd vdd FILL
XFILL_60_DFFSR_255 gnd vdd FILL
XFILL_14_NOR3X1_21 gnd vdd FILL
XFILL_37_DFFSR_97 gnd vdd FILL
XFILL_60_DFFSR_266 gnd vdd FILL
XFILL_77_DFFSR_30 gnd vdd FILL
XFILL_14_NOR3X1_32 gnd vdd FILL
XFILL_77_DFFSR_41 gnd vdd FILL
XFILL_14_NOR3X1_43 gnd vdd FILL
XFILL_64_DFFSR_210 gnd vdd FILL
XFILL_77_DFFSR_52 gnd vdd FILL
XFILL_77_DFFSR_63 gnd vdd FILL
XFILL_7_BUFX4_101 gnd vdd FILL
XFILL_64_DFFSR_221 gnd vdd FILL
XFILL_38_5_0 gnd vdd FILL
XFILL_77_DFFSR_74 gnd vdd FILL
XFILL_64_DFFSR_232 gnd vdd FILL
XFILL_64_DFFSR_243 gnd vdd FILL
XFILL_77_DFFSR_85 gnd vdd FILL
XFILL_64_DFFSR_254 gnd vdd FILL
XFILL_77_DFFSR_96 gnd vdd FILL
XFILL_18_NOR3X1_20 gnd vdd FILL
XFILL_64_DFFSR_265 gnd vdd FILL
XFILL_4_CLKBUF1_30 gnd vdd FILL
XFILL_18_NOR3X1_31 gnd vdd FILL
XFILL_4_CLKBUF1_41 gnd vdd FILL
XFILL_18_NOR3X1_42 gnd vdd FILL
XFILL_12_MUX2X1_104 gnd vdd FILL
XFILL_0_INVX1_70 gnd vdd FILL
XFILL_12_MUX2X1_115 gnd vdd FILL
XFILL_68_DFFSR_220 gnd vdd FILL
XFILL_0_INVX1_81 gnd vdd FILL
XFILL_12_MUX2X1_126 gnd vdd FILL
XFILL_0_INVX1_92 gnd vdd FILL
XFILL_12_MUX2X1_137 gnd vdd FILL
XFILL_68_DFFSR_231 gnd vdd FILL
XFILL_52_0_2 gnd vdd FILL
XFILL_46_DFFSR_40 gnd vdd FILL
XFILL_68_DFFSR_242 gnd vdd FILL
XFILL_17_NOR3X1_4 gnd vdd FILL
XFILL_46_DFFSR_51 gnd vdd FILL
XFILL_12_MUX2X1_148 gnd vdd FILL
XFILL_68_DFFSR_253 gnd vdd FILL
XFILL_12_MUX2X1_159 gnd vdd FILL
XFILL_68_DFFSR_264 gnd vdd FILL
XFILL_46_DFFSR_62 gnd vdd FILL
XFILL_23_CLKBUF1_5 gnd vdd FILL
XFILL_68_DFFSR_275 gnd vdd FILL
XFILL_46_DFFSR_73 gnd vdd FILL
XFILL_46_DFFSR_84 gnd vdd FILL
XFILL_46_DFFSR_95 gnd vdd FILL
XFILL_1_NOR2X1_15 gnd vdd FILL
XFILL_1_NOR2X1_26 gnd vdd FILL
XFILL_13_OAI21X1_20 gnd vdd FILL
XFILL_1_NOR2X1_37 gnd vdd FILL
XFILL_13_OAI21X1_31 gnd vdd FILL
XFILL_21_4_0 gnd vdd FILL
XFILL_13_OAI21X1_42 gnd vdd FILL
XFILL_1_NOR2X1_48 gnd vdd FILL
XFILL_1_NOR2X1_59 gnd vdd FILL
XFILL_86_DFFSR_50 gnd vdd FILL
XFILL_86_DFFSR_61 gnd vdd FILL
XFILL_27_CLKBUF1_4 gnd vdd FILL
XFILL_2_NOR2X1_170 gnd vdd FILL
XFILL_2_NOR2X1_181 gnd vdd FILL
XFILL_86_DFFSR_72 gnd vdd FILL
XFILL_86_DFFSR_83 gnd vdd FILL
XFILL_2_NOR2X1_192 gnd vdd FILL
XFILL_86_DFFSR_94 gnd vdd FILL
XFILL_5_NOR2X1_14 gnd vdd FILL
XFILL_15_DFFSR_50 gnd vdd FILL
XFILL_5_NOR2X1_25 gnd vdd FILL
XFILL_15_DFFSR_61 gnd vdd FILL
XFILL_5_NOR2X1_36 gnd vdd FILL
XFILL_5_NOR2X1_47 gnd vdd FILL
XFILL_15_DFFSR_72 gnd vdd FILL
XFILL_15_DFFSR_83 gnd vdd FILL
XFILL_5_NOR2X1_58 gnd vdd FILL
XFILL_15_DFFSR_94 gnd vdd FILL
XFILL_5_NOR2X1_69 gnd vdd FILL
XFILL_26_NOR3X1_2 gnd vdd FILL
XFILL_9_NOR2X1_13 gnd vdd FILL
XFILL_55_DFFSR_60 gnd vdd FILL
XFILL_9_NOR2X1_24 gnd vdd FILL
XFILL_9_NOR2X1_35 gnd vdd FILL
XFILL_55_DFFSR_71 gnd vdd FILL
XFILL_9_NOR2X1_46 gnd vdd FILL
XFILL_55_DFFSR_82 gnd vdd FILL
XFILL_9_NOR2X1_57 gnd vdd FILL
XFILL_13_OAI22X1_8 gnd vdd FILL
XFILL_55_DFFSR_93 gnd vdd FILL
XFILL_9_NOR2X1_68 gnd vdd FILL
XFILL_9_NOR2X1_79 gnd vdd FILL
XFILL_2_MUX2X1_110 gnd vdd FILL
XFILL_0_NOR2X1_3 gnd vdd FILL
XFILL_2_MUX2X1_121 gnd vdd FILL
XFILL_77_DFFSR_109 gnd vdd FILL
XFILL_2_MUX2X1_132 gnd vdd FILL
XFILL_2_MUX2X1_143 gnd vdd FILL
XFILL_2_MUX2X1_154 gnd vdd FILL
XFILL_2_MUX2X1_165 gnd vdd FILL
XFILL_17_OAI22X1_7 gnd vdd FILL
XFILL_15_NAND3X1_18 gnd vdd FILL
XFILL_15_NAND3X1_29 gnd vdd FILL
XFILL_2_MUX2X1_176 gnd vdd FILL
XFILL_2_MUX2X1_187 gnd vdd FILL
XFILL_24_DFFSR_70 gnd vdd FILL
XFILL_24_DFFSR_81 gnd vdd FILL
XFILL_29_5_0 gnd vdd FILL
XFILL_24_DFFSR_92 gnd vdd FILL
XFILL_4_5_0 gnd vdd FILL
XFILL_9_NOR3X1_3 gnd vdd FILL
XFILL_35_CLKBUF1_18 gnd vdd FILL
XFILL_31_DFFSR_210 gnd vdd FILL
XFILL_35_CLKBUF1_29 gnd vdd FILL
XFILL_7_BUFX2_3 gnd vdd FILL
XFILL_31_DFFSR_221 gnd vdd FILL
XFILL_31_DFFSR_232 gnd vdd FILL
XFILL_31_DFFSR_243 gnd vdd FILL
XFILL_31_DFFSR_254 gnd vdd FILL
XFILL_64_DFFSR_80 gnd vdd FILL
XFILL_31_DFFSR_265 gnd vdd FILL
XFILL_64_DFFSR_91 gnd vdd FILL
XFILL_43_0_2 gnd vdd FILL
XFILL_35_DFFSR_220 gnd vdd FILL
XFILL_35_DFFSR_231 gnd vdd FILL
XFILL_35_DFFSR_242 gnd vdd FILL
XFILL_35_DFFSR_253 gnd vdd FILL
XFILL_66_DFFSR_2 gnd vdd FILL
XFILL_35_DFFSR_264 gnd vdd FILL
XFILL_7_DFFSR_60 gnd vdd FILL
XFILL_1_MUX2X1_11 gnd vdd FILL
XFILL_35_DFFSR_275 gnd vdd FILL
XFILL_1_MUX2X1_22 gnd vdd FILL
XFILL_12_4_0 gnd vdd FILL
XFILL_7_DFFSR_71 gnd vdd FILL
XFILL_7_DFFSR_82 gnd vdd FILL
XFILL_1_MUX2X1_33 gnd vdd FILL
XINVX8_1 din[1] gnd INVX8_1/Y vdd INVX8
XFILL_1_MUX2X1_44 gnd vdd FILL
XFILL_7_DFFSR_93 gnd vdd FILL
XFILL_62_DFFSR_120 gnd vdd FILL
XFILL_62_DFFSR_131 gnd vdd FILL
XFILL_1_MUX2X1_55 gnd vdd FILL
XFILL_33_DFFSR_90 gnd vdd FILL
XFILL_62_DFFSR_142 gnd vdd FILL
XFILL_1_MUX2X1_66 gnd vdd FILL
XFILL_39_DFFSR_230 gnd vdd FILL
XFILL_1_MUX2X1_77 gnd vdd FILL
XFILL_39_DFFSR_241 gnd vdd FILL
XFILL_1_MUX2X1_88 gnd vdd FILL
XFILL_62_DFFSR_153 gnd vdd FILL
XFILL_39_DFFSR_252 gnd vdd FILL
XFILL_14_NAND3X1_109 gnd vdd FILL
XFILL_39_DFFSR_263 gnd vdd FILL
XFILL_62_DFFSR_164 gnd vdd FILL
XFILL_39_DFFSR_274 gnd vdd FILL
XFILL_1_MUX2X1_99 gnd vdd FILL
XFILL_62_DFFSR_175 gnd vdd FILL
XFILL_5_MUX2X1_10 gnd vdd FILL
XFILL_5_MUX2X1_21 gnd vdd FILL
XFILL_62_DFFSR_186 gnd vdd FILL
XFILL_62_DFFSR_197 gnd vdd FILL
XFILL_5_MUX2X1_32 gnd vdd FILL
XFILL_5_MUX2X1_43 gnd vdd FILL
XFILL_5_MUX2X1_54 gnd vdd FILL
XFILL_5_NAND3X1_13 gnd vdd FILL
XFILL_66_DFFSR_130 gnd vdd FILL
XFILL_5_NAND3X1_24 gnd vdd FILL
XFILL_5_MUX2X1_65 gnd vdd FILL
XFILL_5_NAND3X1_35 gnd vdd FILL
XFILL_66_DFFSR_141 gnd vdd FILL
XFILL_66_DFFSR_152 gnd vdd FILL
XFILL_5_MUX2X1_76 gnd vdd FILL
XFILL_5_MUX2X1_87 gnd vdd FILL
XFILL_5_NAND3X1_46 gnd vdd FILL
XFILL_5_NAND3X1_57 gnd vdd FILL
XFILL_50_DFFSR_8 gnd vdd FILL
XFILL_66_DFFSR_163 gnd vdd FILL
XFILL_5_MUX2X1_98 gnd vdd FILL
XFILL_9_NAND2X1_15 gnd vdd FILL
XFILL_66_DFFSR_174 gnd vdd FILL
XFILL_5_NAND3X1_68 gnd vdd FILL
XFILL_9_NAND2X1_26 gnd vdd FILL
XFILL_5_NAND3X1_79 gnd vdd FILL
XFILL_9_MUX2X1_20 gnd vdd FILL
XFILL_66_DFFSR_185 gnd vdd FILL
XFILL_9_MUX2X1_31 gnd vdd FILL
XFILL_9_NAND2X1_37 gnd vdd FILL
XFILL_66_DFFSR_196 gnd vdd FILL
XFILL_9_NAND2X1_48 gnd vdd FILL
XFILL_9_MUX2X1_42 gnd vdd FILL
XFILL_17_DFFSR_209 gnd vdd FILL
XFILL_9_MUX2X1_53 gnd vdd FILL
XFILL_9_NAND2X1_59 gnd vdd FILL
XFILL_14_NAND3X1_9 gnd vdd FILL
XFILL_9_MUX2X1_64 gnd vdd FILL
XFILL_9_MUX2X1_75 gnd vdd FILL
XFILL_9_MUX2X1_86 gnd vdd FILL
XFILL_9_MUX2X1_97 gnd vdd FILL
XFILL_7_INVX2_3 gnd vdd FILL
XBUFX4_10 clk gnd BUFX4_10/Y vdd BUFX4
XFILL_44_DFFSR_109 gnd vdd FILL
XBUFX4_21 BUFX4_51/Y gnd BUFX4_21/Y vdd BUFX4
XFILL_19_MUX2X1_190 gnd vdd FILL
XBUFX4_32 BUFX4_44/A gnd BUFX4_32/Y vdd BUFX4
XBUFX4_43 BUFX4_3/Y gnd DFFSR_73/R vdd BUFX4
XBUFX4_54 BUFX4_54/A gnd BUFX4_54/Y vdd BUFX4
XBUFX4_65 INVX8_1/Y gnd BUFX4_65/Y vdd BUFX4
XBUFX4_76 INVX8_2/Y gnd BUFX4_76/Y vdd BUFX4
XBUFX4_87 INVX8_4/Y gnd BUFX4_87/Y vdd BUFX4
XBUFX4_98 INVX8_3/Y gnd BUFX4_98/Y vdd BUFX4
XFILL_48_DFFSR_108 gnd vdd FILL
XFILL_5_INVX1_1 gnd vdd FILL
XFILL_21_MUX2X1_30 gnd vdd FILL
XFILL_48_DFFSR_119 gnd vdd FILL
XFILL_21_MUX2X1_41 gnd vdd FILL
XFILL_21_MUX2X1_52 gnd vdd FILL
XFILL_62_3_0 gnd vdd FILL
XFILL_21_MUX2X1_63 gnd vdd FILL
XFILL_34_0_2 gnd vdd FILL
XFILL_21_MUX2X1_74 gnd vdd FILL
XFILL_21_MUX2X1_85 gnd vdd FILL
XFILL_21_MUX2X1_96 gnd vdd FILL
XFILL_10_2 gnd vdd FILL
XFILL_24_CLKBUF1_14 gnd vdd FILL
XFILL_24_CLKBUF1_25 gnd vdd FILL
XFILL_24_CLKBUF1_36 gnd vdd FILL
XFILL_7_CLKBUF1_18 gnd vdd FILL
XFILL_7_CLKBUF1_29 gnd vdd FILL
XFILL_10_AND2X2_8 gnd vdd FILL
XFILL_33_DFFSR_130 gnd vdd FILL
XFILL_2_AOI21X1_15 gnd vdd FILL
XFILL_2_AOI21X1_26 gnd vdd FILL
XFILL_33_DFFSR_141 gnd vdd FILL
XFILL_2_AOI21X1_37 gnd vdd FILL
XFILL_33_DFFSR_152 gnd vdd FILL
XFILL_2_AOI21X1_48 gnd vdd FILL
XFILL_2_AOI21X1_59 gnd vdd FILL
XFILL_33_DFFSR_163 gnd vdd FILL
XFILL_33_DFFSR_174 gnd vdd FILL
XFILL_12_OAI22X1_17 gnd vdd FILL
XFILL_12_OAI22X1_28 gnd vdd FILL
XFILL_33_DFFSR_185 gnd vdd FILL
XFILL_12_OAI22X1_39 gnd vdd FILL
XFILL_33_DFFSR_196 gnd vdd FILL
XFILL_5_NOR2X1_103 gnd vdd FILL
XFILL_5_NOR2X1_114 gnd vdd FILL
XFILL_5_NOR2X1_125 gnd vdd FILL
XFILL_37_DFFSR_140 gnd vdd FILL
XFILL_37_DFFSR_151 gnd vdd FILL
XFILL_5_NOR2X1_136 gnd vdd FILL
XFILL_5_NOR2X1_147 gnd vdd FILL
XFILL_37_DFFSR_162 gnd vdd FILL
XFILL_5_NOR2X1_158 gnd vdd FILL
XFILL_37_DFFSR_173 gnd vdd FILL
XFILL_37_DFFSR_184 gnd vdd FILL
XFILL_5_NOR2X1_169 gnd vdd FILL
XFILL_11_NAND3X1_60 gnd vdd FILL
XFILL_37_DFFSR_195 gnd vdd FILL
XFILL_11_DFFSR_109 gnd vdd FILL
XFILL_11_NAND3X1_71 gnd vdd FILL
XFILL_11_NAND3X1_82 gnd vdd FILL
XFILL_11_NAND3X1_93 gnd vdd FILL
XFILL_15_DFFSR_108 gnd vdd FILL
XFILL_53_3_0 gnd vdd FILL
XFILL_15_DFFSR_119 gnd vdd FILL
XFILL_25_0_2 gnd vdd FILL
XFILL_0_0_2 gnd vdd FILL
XFILL_22_MUX2X1_105 gnd vdd FILL
XFILL_22_MUX2X1_116 gnd vdd FILL
XFILL_78_DFFSR_19 gnd vdd FILL
XFILL_22_MUX2X1_127 gnd vdd FILL
XFILL_10_DFFSR_1 gnd vdd FILL
XFILL_22_MUX2X1_138 gnd vdd FILL
XFILL_83_DFFSR_230 gnd vdd FILL
XFILL_10_AOI21X1_4 gnd vdd FILL
XFILL_22_MUX2X1_149 gnd vdd FILL
XFILL_83_DFFSR_241 gnd vdd FILL
XFILL_83_DFFSR_252 gnd vdd FILL
XFILL_83_DFFSR_263 gnd vdd FILL
XFILL_5_MUX2X1_109 gnd vdd FILL
XFILL_83_DFFSR_274 gnd vdd FILL
XFILL_19_DFFSR_107 gnd vdd FILL
XFILL_19_DFFSR_118 gnd vdd FILL
XFILL_1_INVX1_15 gnd vdd FILL
XFILL_19_DFFSR_129 gnd vdd FILL
XFILL_1_INVX1_26 gnd vdd FILL
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XFILL_1_INVX1_37 gnd vdd FILL
XFILL_14_AOI21X1_3 gnd vdd FILL
XFILL_2_OAI22X1_12 gnd vdd FILL
XFILL_1_INVX1_48 gnd vdd FILL
XFILL_2_AND2X2_7 gnd vdd FILL
XFILL_1_INVX1_59 gnd vdd FILL
XFILL_2_OAI22X1_23 gnd vdd FILL
XFILL_87_DFFSR_240 gnd vdd FILL
XFILL_87_DFFSR_251 gnd vdd FILL
XFILL_2_OAI22X1_34 gnd vdd FILL
XFILL_87_DFFSR_262 gnd vdd FILL
XFILL_2_OAI22X1_45 gnd vdd FILL
XFILL_87_DFFSR_273 gnd vdd FILL
XFILL_47_DFFSR_18 gnd vdd FILL
XFILL_6_OAI21X1_14 gnd vdd FILL
XFILL_47_DFFSR_29 gnd vdd FILL
XFILL_6_OAI21X1_25 gnd vdd FILL
XFILL_6_OAI21X1_36 gnd vdd FILL
XFILL_6_OAI21X1_47 gnd vdd FILL
XFILL_61_DFFSR_209 gnd vdd FILL
XFILL_3_INVX1_190 gnd vdd FILL
XFILL_15_NOR3X1_19 gnd vdd FILL
XFILL_87_DFFSR_17 gnd vdd FILL
XFILL_87_DFFSR_28 gnd vdd FILL
XFILL_32_DFFSR_5 gnd vdd FILL
XFILL_87_DFFSR_39 gnd vdd FILL
XFILL_65_DFFSR_208 gnd vdd FILL
XFILL_65_DFFSR_219 gnd vdd FILL
XFILL_16_DFFSR_17 gnd vdd FILL
XFILL_16_DFFSR_28 gnd vdd FILL
XFILL_16_DFFSR_39 gnd vdd FILL
XFILL_5_NAND2X1_90 gnd vdd FILL
XFILL_19_NOR3X1_18 gnd vdd FILL
XFILL_8_1_2 gnd vdd FILL
XFILL_19_NOR3X1_29 gnd vdd FILL
XFILL_13_CLKBUF1_10 gnd vdd FILL
XFILL_69_DFFSR_207 gnd vdd FILL
XFILL_13_CLKBUF1_21 gnd vdd FILL
XFILL_13_CLKBUF1_32 gnd vdd FILL
XFILL_69_DFFSR_218 gnd vdd FILL
XFILL_56_DFFSR_16 gnd vdd FILL
XFILL_56_DFFSR_27 gnd vdd FILL
XFILL_69_DFFSR_229 gnd vdd FILL
XFILL_56_DFFSR_38 gnd vdd FILL
XFILL_56_DFFSR_49 gnd vdd FILL
XFILL_44_3_0 gnd vdd FILL
XFILL_16_0_2 gnd vdd FILL
XFILL_54_DFFSR_9 gnd vdd FILL
XFILL_25_DFFSR_15 gnd vdd FILL
XFILL_11_NOR2X1_150 gnd vdd FILL
XFILL_25_DFFSR_26 gnd vdd FILL
XFILL_11_NOR2X1_161 gnd vdd FILL
XFILL_25_DFFSR_37 gnd vdd FILL
XFILL_25_DFFSR_48 gnd vdd FILL
XFILL_11_NOR2X1_172 gnd vdd FILL
XFILL_11_NOR2X1_183 gnd vdd FILL
XFILL_25_DFFSR_59 gnd vdd FILL
XFILL_11_NOR2X1_194 gnd vdd FILL
XFILL_50_DFFSR_230 gnd vdd FILL
XFILL_50_DFFSR_241 gnd vdd FILL
XFILL_65_DFFSR_14 gnd vdd FILL
XFILL_50_DFFSR_252 gnd vdd FILL
XFILL_65_DFFSR_25 gnd vdd FILL
XFILL_50_DFFSR_263 gnd vdd FILL
XFILL_50_DFFSR_274 gnd vdd FILL
XFILL_65_DFFSR_36 gnd vdd FILL
XFILL_65_DFFSR_47 gnd vdd FILL
XFILL_65_DFFSR_58 gnd vdd FILL
XFILL_65_DFFSR_69 gnd vdd FILL
XFILL_54_DFFSR_240 gnd vdd FILL
XFILL_54_DFFSR_251 gnd vdd FILL
XFILL_54_DFFSR_262 gnd vdd FILL
XFILL_8_DFFSR_16 gnd vdd FILL
XFILL_54_DFFSR_273 gnd vdd FILL
XFILL_8_DFFSR_27 gnd vdd FILL
XFILL_11_MUX2X1_101 gnd vdd FILL
XFILL_34_DFFSR_13 gnd vdd FILL
XFILL_8_DFFSR_38 gnd vdd FILL
XFILL_11_MUX2X1_112 gnd vdd FILL
XFILL_34_DFFSR_24 gnd vdd FILL
XFILL_8_DFFSR_49 gnd vdd FILL
XFILL_11_MUX2X1_123 gnd vdd FILL
XFILL_34_DFFSR_35 gnd vdd FILL
XFILL_81_DFFSR_140 gnd vdd FILL
XFILL_11_MUX2X1_134 gnd vdd FILL
XFILL_11_MUX2X1_145 gnd vdd FILL
XFILL_34_DFFSR_46 gnd vdd FILL
XFILL_34_DFFSR_57 gnd vdd FILL
XFILL_81_DFFSR_151 gnd vdd FILL
XFILL_58_DFFSR_250 gnd vdd FILL
XFILL_81_DFFSR_162 gnd vdd FILL
XFILL_11_MUX2X1_156 gnd vdd FILL
XFILL_34_DFFSR_68 gnd vdd FILL
XFILL_58_DFFSR_261 gnd vdd FILL
XFILL_58_DFFSR_272 gnd vdd FILL
XFILL_81_DFFSR_173 gnd vdd FILL
XFILL_34_DFFSR_79 gnd vdd FILL
XFILL_11_MUX2X1_167 gnd vdd FILL
XFILL_13_CLKBUF1_2 gnd vdd FILL
XFILL_81_DFFSR_184 gnd vdd FILL
XFILL_11_MUX2X1_178 gnd vdd FILL
XFILL_11_MUX2X1_189 gnd vdd FILL
XFILL_1_DFFSR_210 gnd vdd FILL
XFILL_81_DFFSR_195 gnd vdd FILL
XFILL_32_DFFSR_208 gnd vdd FILL
XFILL_74_DFFSR_12 gnd vdd FILL
XFILL_1_DFFSR_221 gnd vdd FILL
XFILL_74_DFFSR_23 gnd vdd FILL
XFILL_32_DFFSR_219 gnd vdd FILL
XFILL_9_1 gnd vdd FILL
XFILL_1_DFFSR_232 gnd vdd FILL
XFILL_74_DFFSR_34 gnd vdd FILL
XFILL_1_DFFSR_243 gnd vdd FILL
XFILL_74_DFFSR_45 gnd vdd FILL
XFILL_17_MUX2X1_2 gnd vdd FILL
XFILL_1_DFFSR_254 gnd vdd FILL
XFILL_85_DFFSR_150 gnd vdd FILL
XFILL_74_DFFSR_56 gnd vdd FILL
XFILL_12_OAI21X1_50 gnd vdd FILL
XFILL_1_DFFSR_265 gnd vdd FILL
XFILL_85_DFFSR_161 gnd vdd FILL
XFILL_74_DFFSR_67 gnd vdd FILL
XFILL_74_DFFSR_78 gnd vdd FILL
XFILL_17_CLKBUF1_1 gnd vdd FILL
XFILL_85_DFFSR_172 gnd vdd FILL
XFILL_65_3 gnd vdd FILL
XFILL_74_DFFSR_89 gnd vdd FILL
XFILL_85_DFFSR_183 gnd vdd FILL
XFILL_85_DFFSR_194 gnd vdd FILL
XFILL_36_DFFSR_207 gnd vdd FILL
XFILL_5_DFFSR_220 gnd vdd FILL
XFILL_36_DFFSR_218 gnd vdd FILL
XFILL_58_2 gnd vdd FILL
XFILL_5_DFFSR_231 gnd vdd FILL
XFILL_5_DFFSR_242 gnd vdd FILL
XFILL_36_DFFSR_229 gnd vdd FILL
XFILL_5_DFFSR_253 gnd vdd FILL
XFILL_43_DFFSR_11 gnd vdd FILL
XFILL_5_DFFSR_264 gnd vdd FILL
XFILL_43_DFFSR_22 gnd vdd FILL
XFILL_5_DFFSR_275 gnd vdd FILL
XFILL_43_DFFSR_33 gnd vdd FILL
XFILL_14_NOR3X1_8 gnd vdd FILL
XFILL_8_BUFX4_90 gnd vdd FILL
XFILL_43_DFFSR_44 gnd vdd FILL
XFILL_43_DFFSR_55 gnd vdd FILL
XFILL_35_3_0 gnd vdd FILL
XFILL_63_DFFSR_107 gnd vdd FILL
XFILL_43_DFFSR_66 gnd vdd FILL
XFILL_63_DFFSR_118 gnd vdd FILL
XFILL_43_DFFSR_77 gnd vdd FILL
XFILL_9_DFFSR_230 gnd vdd FILL
XFILL_63_DFFSR_129 gnd vdd FILL
XFILL_9_DFFSR_241 gnd vdd FILL
XFILL_43_DFFSR_88 gnd vdd FILL
XFILL_43_DFFSR_99 gnd vdd FILL
XFILL_9_DFFSR_252 gnd vdd FILL
XFILL_83_DFFSR_10 gnd vdd FILL
XFILL_10_NAND3X1_106 gnd vdd FILL
XFILL_9_DFFSR_263 gnd vdd FILL
XFILL_9_DFFSR_274 gnd vdd FILL
XFILL_83_DFFSR_21 gnd vdd FILL
XFILL_10_NAND3X1_117 gnd vdd FILL
XFILL_10_NAND3X1_128 gnd vdd FILL
XFILL_83_DFFSR_32 gnd vdd FILL
XFILL_83_DFFSR_43 gnd vdd FILL
XFILL_6_MUX2X1_19 gnd vdd FILL
XFILL_12_DFFSR_10 gnd vdd FILL
XFILL_83_DFFSR_54 gnd vdd FILL
XFILL_67_DFFSR_106 gnd vdd FILL
XFILL_83_DFFSR_65 gnd vdd FILL
XFILL_12_DFFSR_21 gnd vdd FILL
XFILL_67_DFFSR_117 gnd vdd FILL
XFILL_83_DFFSR_76 gnd vdd FILL
XFILL_1_MUX2X1_140 gnd vdd FILL
XFILL_12_DFFSR_32 gnd vdd FILL
XFILL_67_DFFSR_128 gnd vdd FILL
XFILL_12_DFFSR_43 gnd vdd FILL
XFILL_83_DFFSR_87 gnd vdd FILL
XFILL_67_DFFSR_139 gnd vdd FILL
XFILL_1_MUX2X1_151 gnd vdd FILL
XFILL_1_MUX2X1_162 gnd vdd FILL
XFILL_83_DFFSR_98 gnd vdd FILL
XFILL_14_NAND3X1_15 gnd vdd FILL
XFILL_12_DFFSR_54 gnd vdd FILL
XFILL_1_MUX2X1_173 gnd vdd FILL
XFILL_10_OAI21X1_7 gnd vdd FILL
XFILL_12_DFFSR_65 gnd vdd FILL
XFILL_14_NAND3X1_26 gnd vdd FILL
XFILL_12_DFFSR_76 gnd vdd FILL
XFILL_14_NAND3X1_37 gnd vdd FILL
XFILL_1_MUX2X1_184 gnd vdd FILL
XFILL_12_DFFSR_87 gnd vdd FILL
XFILL_14_NAND3X1_48 gnd vdd FILL
XFILL_14_NAND3X1_59 gnd vdd FILL
XFILL_12_DFFSR_98 gnd vdd FILL
XFILL_52_DFFSR_20 gnd vdd FILL
XFILL_34_CLKBUF1_15 gnd vdd FILL
XFILL_34_CLKBUF1_26 gnd vdd FILL
XFILL_52_DFFSR_31 gnd vdd FILL
XFILL_23_NOR3X1_6 gnd vdd FILL
XFILL_52_DFFSR_42 gnd vdd FILL
XFILL_11_NOR2X1_20 gnd vdd FILL
XFILL_2_AOI22X1_3 gnd vdd FILL
XFILL_34_CLKBUF1_37 gnd vdd FILL
XFILL_14_OAI21X1_6 gnd vdd FILL
XFILL_11_NOR2X1_31 gnd vdd FILL
XFILL_52_DFFSR_53 gnd vdd FILL
XFILL_11_NOR2X1_42 gnd vdd FILL
XFILL_21_DFFSR_240 gnd vdd FILL
XFILL_52_DFFSR_64 gnd vdd FILL
XFILL_11_NOR2X1_53 gnd vdd FILL
XFILL_21_DFFSR_251 gnd vdd FILL
XFILL_52_DFFSR_75 gnd vdd FILL
XFILL_21_DFFSR_262 gnd vdd FILL
XFILL_52_DFFSR_86 gnd vdd FILL
XFILL_11_NOR2X1_64 gnd vdd FILL
XFILL_11_NOR2X1_75 gnd vdd FILL
XFILL_2_INVX1_202 gnd vdd FILL
XFILL_21_DFFSR_273 gnd vdd FILL
XFILL_52_DFFSR_97 gnd vdd FILL
XFILL_2_INVX1_213 gnd vdd FILL
XFILL_11_NOR2X1_86 gnd vdd FILL
XFILL_1_DFFSR_4 gnd vdd FILL
XFILL_9_MUX2X1_1 gnd vdd FILL
XFILL_11_NOR2X1_97 gnd vdd FILL
XFILL_2_INVX1_224 gnd vdd FILL
XFILL_6_AOI22X1_2 gnd vdd FILL
XFILL_14_DFFSR_2 gnd vdd FILL
XFILL_71_DFFSR_3 gnd vdd FILL
XFILL_21_DFFSR_30 gnd vdd FILL
XFILL_25_DFFSR_250 gnd vdd FILL
XFILL_25_DFFSR_261 gnd vdd FILL
XFILL_25_DFFSR_272 gnd vdd FILL
XFILL_21_DFFSR_41 gnd vdd FILL
XFILL_21_DFFSR_52 gnd vdd FILL
XFILL_6_INVX1_201 gnd vdd FILL
XFILL_21_DFFSR_63 gnd vdd FILL
XFILL_6_INVX1_212 gnd vdd FILL
XFILL_22_MUX2X1_17 gnd vdd FILL
XFILL_6_INVX1_223 gnd vdd FILL
XFILL_21_DFFSR_74 gnd vdd FILL
XFILL_22_MUX2X1_28 gnd vdd FILL
XFILL_21_DFFSR_85 gnd vdd FILL
XFILL_22_MUX2X1_39 gnd vdd FILL
XFILL_21_DFFSR_96 gnd vdd FILL
XFILL_52_DFFSR_150 gnd vdd FILL
XFILL_6_NOR3X1_7 gnd vdd FILL
XFILL_52_DFFSR_161 gnd vdd FILL
XFILL_61_DFFSR_40 gnd vdd FILL
XFILL_29_DFFSR_260 gnd vdd FILL
XFILL_29_DFFSR_271 gnd vdd FILL
XFILL_52_DFFSR_172 gnd vdd FILL
XFILL_61_DFFSR_51 gnd vdd FILL
XFILL_52_DFFSR_183 gnd vdd FILL
XFILL_52_DFFSR_194 gnd vdd FILL
XFILL_61_DFFSR_62 gnd vdd FILL
XFILL_61_DFFSR_73 gnd vdd FILL
XFILL_61_DFFSR_84 gnd vdd FILL
XFILL_4_NAND3X1_10 gnd vdd FILL
XFILL_61_DFFSR_95 gnd vdd FILL
XFILL_4_NAND3X1_21 gnd vdd FILL
XFILL_4_NAND3X1_32 gnd vdd FILL
XFILL_4_NAND3X1_43 gnd vdd FILL
XFILL_56_DFFSR_160 gnd vdd FILL
XFILL_26_3_0 gnd vdd FILL
XFILL_4_DFFSR_20 gnd vdd FILL
XFILL_1_3_0 gnd vdd FILL
XFILL_8_NAND2X1_12 gnd vdd FILL
XFILL_4_NAND3X1_54 gnd vdd FILL
XFILL_4_NAND3X1_65 gnd vdd FILL
XFILL_8_NAND2X1_23 gnd vdd FILL
XFILL_4_DFFSR_31 gnd vdd FILL
XFILL_56_DFFSR_171 gnd vdd FILL
XFILL_4_NAND3X1_76 gnd vdd FILL
XFILL_56_DFFSR_182 gnd vdd FILL
XFILL_4_NAND3X1_87 gnd vdd FILL
XFILL_36_DFFSR_6 gnd vdd FILL
XFILL_4_DFFSR_42 gnd vdd FILL
XFILL_56_DFFSR_193 gnd vdd FILL
XFILL_8_NAND2X1_34 gnd vdd FILL
XFILL_30_DFFSR_107 gnd vdd FILL
XFILL_4_DFFSR_53 gnd vdd FILL
XFILL_8_NAND2X1_45 gnd vdd FILL
XFILL_30_DFFSR_118 gnd vdd FILL
XFILL_4_DFFSR_64 gnd vdd FILL
XFILL_8_NAND2X1_56 gnd vdd FILL
XFILL_4_NAND3X1_98 gnd vdd FILL
XFILL_4_DFFSR_75 gnd vdd FILL
XFILL_30_DFFSR_129 gnd vdd FILL
XFILL_8_NAND2X1_67 gnd vdd FILL
XFILL_30_DFFSR_50 gnd vdd FILL
XFILL_4_DFFSR_86 gnd vdd FILL
XFILL_8_NAND2X1_78 gnd vdd FILL
XFILL_30_DFFSR_61 gnd vdd FILL
XFILL_8_NAND2X1_89 gnd vdd FILL
XFILL_30_DFFSR_72 gnd vdd FILL
XFILL_4_DFFSR_97 gnd vdd FILL
XFILL_30_DFFSR_83 gnd vdd FILL
XFILL_30_DFFSR_94 gnd vdd FILL
XFILL_34_DFFSR_106 gnd vdd FILL
XFILL_3_DFFSR_130 gnd vdd FILL
XFILL_34_DFFSR_117 gnd vdd FILL
XFILL_11_NAND2X1_8 gnd vdd FILL
XFILL_10_7_1 gnd vdd FILL
XFILL_34_DFFSR_128 gnd vdd FILL
XFILL_3_DFFSR_141 gnd vdd FILL
XFILL_3_DFFSR_152 gnd vdd FILL
XFILL_70_DFFSR_60 gnd vdd FILL
XFILL_34_DFFSR_139 gnd vdd FILL
XFILL_11_AOI21X1_17 gnd vdd FILL
XFILL_3_DFFSR_163 gnd vdd FILL
XFILL_70_DFFSR_71 gnd vdd FILL
XFILL_70_DFFSR_82 gnd vdd FILL
XFILL_3_DFFSR_174 gnd vdd FILL
XFILL_11_AOI21X1_28 gnd vdd FILL
XFILL_70_DFFSR_93 gnd vdd FILL
XFILL_11_AOI21X1_39 gnd vdd FILL
XFILL_3_DFFSR_185 gnd vdd FILL
XFILL_3_DFFSR_196 gnd vdd FILL
XFILL_38_DFFSR_105 gnd vdd FILL
XAND2X2_8 INVX4_1/A AND2X2_8/B gnd MUX2X1_1/S vdd AND2X2
XFILL_38_DFFSR_116 gnd vdd FILL
XFILL_7_DFFSR_140 gnd vdd FILL
XFILL_38_DFFSR_127 gnd vdd FILL
XFILL_38_DFFSR_138 gnd vdd FILL
XFILL_7_DFFSR_151 gnd vdd FILL
XFILL_38_DFFSR_149 gnd vdd FILL
XFILL_7_DFFSR_162 gnd vdd FILL
XFILL_10_NOR3X1_1 gnd vdd FILL
XFILL_11_MUX2X1_60 gnd vdd FILL
XFILL_11_MUX2X1_71 gnd vdd FILL
XFILL_7_DFFSR_173 gnd vdd FILL
XFILL_7_DFFSR_184 gnd vdd FILL
XFILL_11_MUX2X1_82 gnd vdd FILL
XFILL_8_AOI22X1_10 gnd vdd FILL
XFILL_11_MUX2X1_93 gnd vdd FILL
XFILL_30_NOR3X1_18 gnd vdd FILL
XFILL_7_DFFSR_195 gnd vdd FILL
XFILL_30_NOR3X1_29 gnd vdd FILL
XFILL_9_4_0 gnd vdd FILL
XFILL_80_DFFSR_207 gnd vdd FILL
XFILL_80_DFFSR_218 gnd vdd FILL
XFILL_80_DFFSR_229 gnd vdd FILL
XFILL_15_MUX2X1_70 gnd vdd FILL
XFILL_15_MUX2X1_81 gnd vdd FILL
XFILL_15_MUX2X1_92 gnd vdd FILL
XFILL_3_NOR3X1_30 gnd vdd FILL
XFILL_3_NOR3X1_41 gnd vdd FILL
XFILL_23_CLKBUF1_11 gnd vdd FILL
XFILL_3_NOR3X1_52 gnd vdd FILL
XFILL_84_DFFSR_206 gnd vdd FILL
XFILL_23_CLKBUF1_22 gnd vdd FILL
XFILL_84_DFFSR_217 gnd vdd FILL
XFILL_23_CLKBUF1_33 gnd vdd FILL
XFILL_84_DFFSR_228 gnd vdd FILL
XFILL_84_DFFSR_239 gnd vdd FILL
XFILL_19_MUX2X1_80 gnd vdd FILL
XFILL_19_MUX2X1_91 gnd vdd FILL
XFILL_6_CLKBUF1_15 gnd vdd FILL
XFILL_6_CLKBUF1_26 gnd vdd FILL
XFILL_7_NOR3X1_40 gnd vdd FILL
XFILL_0_INVX1_101 gnd vdd FILL
XFILL_0_INVX1_112 gnd vdd FILL
XFILL_0_INVX1_123 gnd vdd FILL
XFILL_7_NOR3X1_51 gnd vdd FILL
XFILL_17_3_0 gnd vdd FILL
XFILL_6_CLKBUF1_37 gnd vdd FILL
XFILL_1_AOI21X1_12 gnd vdd FILL
XFILL_0_INVX1_134 gnd vdd FILL
XFILL_0_INVX1_145 gnd vdd FILL
XFILL_1_AOI21X1_23 gnd vdd FILL
XFILL_1_AOI21X1_34 gnd vdd FILL
XFILL_0_INVX1_156 gnd vdd FILL
XFILL_0_INVX1_167 gnd vdd FILL
XFILL_1_AOI21X1_45 gnd vdd FILL
XFILL_23_DFFSR_160 gnd vdd FILL
XFILL_1_AOI21X1_56 gnd vdd FILL
XFILL_0_INVX1_178 gnd vdd FILL
XFILL_1_AOI21X1_67 gnd vdd FILL
XFILL_4_INVX1_100 gnd vdd FILL
XFILL_0_INVX1_189 gnd vdd FILL
XFILL_11_OAI22X1_14 gnd vdd FILL
XFILL_23_DFFSR_171 gnd vdd FILL
XFILL_60_6_1 gnd vdd FILL
XFILL_11_OAI22X1_25 gnd vdd FILL
XFILL_23_DFFSR_182 gnd vdd FILL
XFILL_1_AOI21X1_78 gnd vdd FILL
XFILL_23_DFFSR_193 gnd vdd FILL
XFILL_11_OAI22X1_36 gnd vdd FILL
XFILL_4_INVX1_111 gnd vdd FILL
XFILL_4_INVX1_122 gnd vdd FILL
XFILL_11_OAI22X1_47 gnd vdd FILL
XFILL_4_NOR2X1_100 gnd vdd FILL
XFILL_4_INVX1_133 gnd vdd FILL
XFILL_4_INVX1_144 gnd vdd FILL
XFILL_15_OAI21X1_16 gnd vdd FILL
XFILL_4_NOR2X1_111 gnd vdd FILL
XFILL_15_OAI21X1_27 gnd vdd FILL
XFILL_4_INVX1_155 gnd vdd FILL
XFILL_4_NOR2X1_122 gnd vdd FILL
XFILL_4_NOR2X1_133 gnd vdd FILL
XFILL_4_NOR2X1_144 gnd vdd FILL
XFILL_15_OAI21X1_38 gnd vdd FILL
XFILL_4_INVX1_166 gnd vdd FILL
XFILL_15_OAI21X1_49 gnd vdd FILL
XFILL_4_NOR2X1_155 gnd vdd FILL
XFILL_4_INVX1_177 gnd vdd FILL
XFILL_4_INVX1_188 gnd vdd FILL
XFILL_27_DFFSR_170 gnd vdd FILL
XFILL_4_INVX1_199 gnd vdd FILL
XFILL_4_NOR2X1_166 gnd vdd FILL
XFILL_27_DFFSR_181 gnd vdd FILL
XFILL_4_NOR2X1_177 gnd vdd FILL
XFILL_27_DFFSR_192 gnd vdd FILL
XFILL_4_NOR2X1_188 gnd vdd FILL
XFILL_4_NOR2X1_199 gnd vdd FILL
XFILL_10_NAND3X1_90 gnd vdd FILL
XFILL_21_MUX2X1_102 gnd vdd FILL
XFILL_21_MUX2X1_113 gnd vdd FILL
XFILL_2_OAI22X1_6 gnd vdd FILL
XFILL_21_MUX2X1_124 gnd vdd FILL
XFILL_21_MUX2X1_135 gnd vdd FILL
XFILL_21_MUX2X1_146 gnd vdd FILL
XFILL_21_MUX2X1_157 gnd vdd FILL
XFILL_73_DFFSR_260 gnd vdd FILL
XFILL_73_DFFSR_271 gnd vdd FILL
XFILL_4_MUX2X1_106 gnd vdd FILL
XFILL_21_MUX2X1_168 gnd vdd FILL
XFILL_4_MUX2X1_117 gnd vdd FILL
XFILL_21_MUX2X1_179 gnd vdd FILL
XFILL_0_DFFSR_90 gnd vdd FILL
XFILL_4_MUX2X1_128 gnd vdd FILL
XFILL_9_NOR2X1_200 gnd vdd FILL
XFILL_4_MUX2X1_139 gnd vdd FILL
XFILL_6_OAI22X1_5 gnd vdd FILL
XFILL_1_OAI22X1_20 gnd vdd FILL
XFILL_1_OAI22X1_31 gnd vdd FILL
XFILL_1_OAI22X1_42 gnd vdd FILL
XFILL_77_DFFSR_270 gnd vdd FILL
XFILL_5_OAI21X1_11 gnd vdd FILL
XFILL_5_OAI21X1_22 gnd vdd FILL
XFILL_51_DFFSR_206 gnd vdd FILL
XFILL_5_OAI21X1_33 gnd vdd FILL
XFILL_5_OAI21X1_44 gnd vdd FILL
XFILL_51_DFFSR_217 gnd vdd FILL
XFILL_51_DFFSR_228 gnd vdd FILL
XFILL_51_DFFSR_239 gnd vdd FILL
XFILL_5_DFFSR_5 gnd vdd FILL
XFILL_55_DFFSR_205 gnd vdd FILL
XFILL_18_DFFSR_3 gnd vdd FILL
XFILL_55_DFFSR_216 gnd vdd FILL
XFILL_51_6_1 gnd vdd FILL
XFILL_55_DFFSR_227 gnd vdd FILL
XFILL_75_DFFSR_4 gnd vdd FILL
XFILL_11_NAND3X1_107 gnd vdd FILL
XFILL_55_DFFSR_238 gnd vdd FILL
XFILL_9_BUFX4_13 gnd vdd FILL
XFILL_50_1_0 gnd vdd FILL
XFILL_55_DFFSR_249 gnd vdd FILL
XFILL_11_NAND3X1_118 gnd vdd FILL
XFILL_9_BUFX4_24 gnd vdd FILL
XFILL_11_NAND3X1_129 gnd vdd FILL
XFILL_9_BUFX4_35 gnd vdd FILL
XFILL_9_BUFX4_46 gnd vdd FILL
XFILL_9_BUFX4_57 gnd vdd FILL
XFILL_82_DFFSR_105 gnd vdd FILL
XFILL_59_DFFSR_204 gnd vdd FILL
XFILL_59_DFFSR_215 gnd vdd FILL
XFILL_9_BUFX4_68 gnd vdd FILL
XFILL_82_DFFSR_116 gnd vdd FILL
XFILL_82_DFFSR_127 gnd vdd FILL
XFILL_59_DFFSR_226 gnd vdd FILL
XFILL_12_CLKBUF1_40 gnd vdd FILL
XFILL_9_BUFX4_79 gnd vdd FILL
XFILL_82_DFFSR_138 gnd vdd FILL
XFILL_82_DFFSR_149 gnd vdd FILL
XFILL_59_DFFSR_237 gnd vdd FILL
XFILL_59_DFFSR_248 gnd vdd FILL
XFILL_59_DFFSR_259 gnd vdd FILL
XFILL_86_DFFSR_104 gnd vdd FILL
XFILL_2_DFFSR_208 gnd vdd FILL
XFILL_2_DFFSR_219 gnd vdd FILL
XFILL_86_DFFSR_115 gnd vdd FILL
XFILL_86_DFFSR_126 gnd vdd FILL
XFILL_86_DFFSR_137 gnd vdd FILL
XFILL_86_DFFSR_148 gnd vdd FILL
XFILL_86_DFFSR_159 gnd vdd FILL
XFILL_6_DFFSR_207 gnd vdd FILL
XFILL_3_NAND3X1_7 gnd vdd FILL
XFILL_6_DFFSR_218 gnd vdd FILL
XFILL_10_NOR2X1_180 gnd vdd FILL
XFILL_10_NOR2X1_191 gnd vdd FILL
XFILL_6_DFFSR_229 gnd vdd FILL
XFILL_14_BUFX4_105 gnd vdd FILL
XFILL_40_DFFSR_260 gnd vdd FILL
XFILL_59_7_1 gnd vdd FILL
XFILL_40_DFFSR_271 gnd vdd FILL
XFILL_7_NAND3X1_6 gnd vdd FILL
XFILL_58_2_0 gnd vdd FILL
XFILL_44_DFFSR_270 gnd vdd FILL
XFILL_12_BUFX4_3 gnd vdd FILL
XFILL_22_DFFSR_19 gnd vdd FILL
XFILL_13_BUFX4_40 gnd vdd FILL
XFILL_13_BUFX4_51 gnd vdd FILL
XFILL_10_MUX2X1_120 gnd vdd FILL
XFILL_13_BUFX4_62 gnd vdd FILL
XFILL_13_BUFX4_73 gnd vdd FILL
XFILL_10_MUX2X1_131 gnd vdd FILL
XFILL_13_BUFX4_84 gnd vdd FILL
XFILL_10_MUX2X1_142 gnd vdd FILL
XFILL_10_MUX2X1_153 gnd vdd FILL
XFILL_13_BUFX4_95 gnd vdd FILL
XFILL_71_DFFSR_170 gnd vdd FILL
XFILL_10_MUX2X1_164 gnd vdd FILL
XFILL_42_6_1 gnd vdd FILL
XFILL_10_MUX2X1_175 gnd vdd FILL
XFILL_71_DFFSR_181 gnd vdd FILL
XFILL_10_MUX2X1_186 gnd vdd FILL
XFILL_62_DFFSR_18 gnd vdd FILL
XFILL_71_DFFSR_192 gnd vdd FILL
XFILL_22_DFFSR_205 gnd vdd FILL
XFILL_41_1_0 gnd vdd FILL
XFILL_62_DFFSR_29 gnd vdd FILL
XFILL_22_DFFSR_216 gnd vdd FILL
XFILL_22_DFFSR_227 gnd vdd FILL
XFILL_22_DFFSR_238 gnd vdd FILL
XFILL_22_DFFSR_249 gnd vdd FILL
XFILL_75_DFFSR_180 gnd vdd FILL
XFILL_75_DFFSR_191 gnd vdd FILL
XFILL_26_DFFSR_204 gnd vdd FILL
XFILL_26_DFFSR_215 gnd vdd FILL
XAOI22X1_3 AOI22X1_3/A AOI22X1_3/B AOI22X1_3/C AOI22X1_3/D gnd NOR3X1_9/A vdd AOI22X1
XFILL_26_DFFSR_226 gnd vdd FILL
XFILL_26_DFFSR_237 gnd vdd FILL
XFILL_31_DFFSR_17 gnd vdd FILL
XFILL_26_DFFSR_248 gnd vdd FILL
XFILL_31_DFFSR_28 gnd vdd FILL
XFILL_31_DFFSR_39 gnd vdd FILL
XFILL_7_INVX1_30 gnd vdd FILL
XFILL_26_DFFSR_259 gnd vdd FILL
XINVX1_202 DFFSR_86/Q gnd INVX1_202/Y vdd INVX1
XINVX1_213 DFFSR_74/Q gnd INVX1_213/Y vdd INVX1
XFILL_7_INVX1_41 gnd vdd FILL
XFILL_79_DFFSR_190 gnd vdd FILL
XFILL_7_INVX1_52 gnd vdd FILL
XINVX1_224 DFFSR_59/Q gnd INVX1_224/Y vdd INVX1
XFILL_53_DFFSR_104 gnd vdd FILL
XFILL_7_INVX1_63 gnd vdd FILL
XFILL_53_DFFSR_115 gnd vdd FILL
XFILL_7_INVX1_74 gnd vdd FILL
XFILL_7_INVX1_85 gnd vdd FILL
XFILL_53_DFFSR_126 gnd vdd FILL
XFILL_53_DFFSR_137 gnd vdd FILL
XFILL_53_DFFSR_148 gnd vdd FILL
XFILL_7_INVX1_96 gnd vdd FILL
XFILL_71_DFFSR_16 gnd vdd FILL
XFILL_71_DFFSR_27 gnd vdd FILL
XFILL_71_DFFSR_38 gnd vdd FILL
XFILL_53_DFFSR_159 gnd vdd FILL
XFILL_71_DFFSR_49 gnd vdd FILL
XFILL_14_MUX2X1_6 gnd vdd FILL
XFILL_57_DFFSR_103 gnd vdd FILL
XFILL_57_DFFSR_114 gnd vdd FILL
XFILL_57_DFFSR_125 gnd vdd FILL
XFILL_57_DFFSR_136 gnd vdd FILL
XFILL_13_NAND3X1_12 gnd vdd FILL
XFILL_57_DFFSR_147 gnd vdd FILL
XNAND2X1_13 INVX1_166/A INVX2_1/A gnd MUX2X1_91/S vdd NAND2X1
XFILL_57_DFFSR_158 gnd vdd FILL
XFILL_0_MUX2X1_170 gnd vdd FILL
XFILL_13_NAND3X1_23 gnd vdd FILL
XFILL_49_2_0 gnd vdd FILL
XNAND2X1_24 BUFX4_6/Y NOR2X1_38/Y gnd OAI22X1_36/B vdd NAND2X1
XFILL_0_MUX2X1_181 gnd vdd FILL
XFILL_5_BUFX4_50 gnd vdd FILL
XFILL_57_DFFSR_169 gnd vdd FILL
XFILL_13_NAND3X1_34 gnd vdd FILL
XNAND2X1_35 BUFX4_104/Y NOR2X1_34/Y gnd OAI22X1_49/B vdd NAND2X1
XFILL_5_BUFX4_61 gnd vdd FILL
XFILL_13_NAND3X1_45 gnd vdd FILL
XFILL_0_MUX2X1_192 gnd vdd FILL
XNAND2X1_46 AND2X2_2/B AND2X2_2/A gnd NOR3X1_5/B vdd NAND2X1
XFILL_2_INVX8_3 gnd vdd FILL
XFILL_0_DFFSR_107 gnd vdd FILL
XNAND2X1_57 BUFX4_104/Y NOR3X1_9/Y gnd OAI21X1_5/B vdd NAND2X1
XFILL_13_NAND3X1_56 gnd vdd FILL
XFILL_5_BUFX4_72 gnd vdd FILL
XFILL_40_DFFSR_15 gnd vdd FILL
XFILL_33_CLKBUF1_12 gnd vdd FILL
XFILL_15_INVX8_1 gnd vdd FILL
XFILL_40_DFFSR_26 gnd vdd FILL
XFILL_0_DFFSR_118 gnd vdd FILL
XFILL_13_NAND3X1_67 gnd vdd FILL
XNAND2X1_68 NAND2X1_68/A NAND2X1_68/B gnd NOR3X1_31/B vdd NAND2X1
XFILL_5_BUFX4_83 gnd vdd FILL
XFILL_40_DFFSR_37 gnd vdd FILL
XFILL_0_DFFSR_129 gnd vdd FILL
XFILL_13_NAND3X1_78 gnd vdd FILL
XNAND2X1_79 INVX1_99/A INVX1_126/Y gnd NAND3X1_18/A vdd NAND2X1
XFILL_33_CLKBUF1_23 gnd vdd FILL
XFILL_40_DFFSR_48 gnd vdd FILL
XFILL_5_BUFX4_94 gnd vdd FILL
XFILL_33_CLKBUF1_34 gnd vdd FILL
XFILL_13_NAND3X1_89 gnd vdd FILL
XFILL_40_DFFSR_59 gnd vdd FILL
XFILL_42_5 gnd vdd FILL
XFILL_11_DFFSR_270 gnd vdd FILL
XFILL_80_DFFSR_14 gnd vdd FILL
XFILL_4_DFFSR_106 gnd vdd FILL
XFILL_4_DFFSR_117 gnd vdd FILL
XFILL_80_DFFSR_25 gnd vdd FILL
XFILL_80_DFFSR_36 gnd vdd FILL
XFILL_4_DFFSR_128 gnd vdd FILL
XFILL_4_DFFSR_139 gnd vdd FILL
XFILL_80_DFFSR_47 gnd vdd FILL
XFILL_80_DFFSR_58 gnd vdd FILL
XFILL_23_MUX2X1_4 gnd vdd FILL
XFILL_80_DFFSR_69 gnd vdd FILL
XFILL_33_6_1 gnd vdd FILL
XFILL_28_3 gnd vdd FILL
XFILL_32_1_0 gnd vdd FILL
XFILL_8_DFFSR_105 gnd vdd FILL
XFILL_57_DFFSR_1 gnd vdd FILL
XFILL_7_NOR2X1_7 gnd vdd FILL
XFILL_8_DFFSR_116 gnd vdd FILL
XFILL_12_MUX2X1_14 gnd vdd FILL
XFILL_12_MUX2X1_25 gnd vdd FILL
XFILL_8_DFFSR_127 gnd vdd FILL
XFILL_8_DFFSR_138 gnd vdd FILL
XFILL_12_MUX2X1_36 gnd vdd FILL
XFILL_8_DFFSR_149 gnd vdd FILL
XFILL_12_MUX2X1_47 gnd vdd FILL
XFILL_3_AOI21X1_1 gnd vdd FILL
XFILL_4_OAI22X1_19 gnd vdd FILL
XFILL_12_MUX2X1_58 gnd vdd FILL
XFILL_12_MUX2X1_69 gnd vdd FILL
XAOI22X1_11 INVX1_132/Y INVX1_130/A INVX1_131/A INVX1_133/Y gnd OAI21X1_48/A vdd AOI22X1
XFILL_11_BUFX2_10 gnd vdd FILL
XFILL_0_NOR3X1_18 gnd vdd FILL
XFILL_42_DFFSR_180 gnd vdd FILL
XFILL_16_MUX2X1_13 gnd vdd FILL
XFILL_0_NOR3X1_29 gnd vdd FILL
XFILL_42_DFFSR_191 gnd vdd FILL
XFILL_16_MUX2X1_24 gnd vdd FILL
XFILL_16_MUX2X1_35 gnd vdd FILL
XFILL_16_MUX2X1_46 gnd vdd FILL
XFILL_16_MUX2X1_57 gnd vdd FILL
XFILL_6_MUX2X1_5 gnd vdd FILL
XNOR3X1_1 NOR3X1_1/A NOR3X1_1/B INVX2_2/Y gnd NOR3X1_1/Y vdd NOR3X1
XFILL_3_NAND3X1_40 gnd vdd FILL
XFILL_16_MUX2X1_68 gnd vdd FILL
XFILL_3_NAND3X1_51 gnd vdd FILL
XFILL_16_MUX2X1_79 gnd vdd FILL
XFILL_4_NOR3X1_17 gnd vdd FILL
XFILL_3_NAND3X1_62 gnd vdd FILL
XFILL_4_NOR3X1_28 gnd vdd FILL
XFILL_7_NAND2X1_20 gnd vdd FILL
XFILL_3_NAND3X1_73 gnd vdd FILL
XFILL_41_DFFSR_7 gnd vdd FILL
XFILL_7_NAND2X1_31 gnd vdd FILL
XFILL_3_NAND3X1_84 gnd vdd FILL
XFILL_46_DFFSR_190 gnd vdd FILL
XFILL_9_DFFSR_6 gnd vdd FILL
XFILL_4_NOR3X1_39 gnd vdd FILL
XFILL_20_DFFSR_104 gnd vdd FILL
XFILL_3_NAND3X1_95 gnd vdd FILL
XFILL_7_NAND2X1_42 gnd vdd FILL
XFILL_7_NAND2X1_53 gnd vdd FILL
XFILL_20_DFFSR_115 gnd vdd FILL
XFILL_20_DFFSR_126 gnd vdd FILL
XFILL_7_NAND2X1_64 gnd vdd FILL
XFILL_20_DFFSR_137 gnd vdd FILL
XFILL_7_NAND2X1_75 gnd vdd FILL
XFILL_79_DFFSR_5 gnd vdd FILL
XFILL_20_DFFSR_148 gnd vdd FILL
XFILL_7_NAND2X1_86 gnd vdd FILL
XFILL_8_NOR3X1_16 gnd vdd FILL
XFILL_20_DFFSR_159 gnd vdd FILL
XFILL_8_NOR3X1_27 gnd vdd FILL
XFILL_8_NOR3X1_38 gnd vdd FILL
XFILL_24_DFFSR_103 gnd vdd FILL
XFILL_8_NOR3X1_49 gnd vdd FILL
XFILL_24_DFFSR_114 gnd vdd FILL
XFILL_15_CLKBUF1_17 gnd vdd FILL
XFILL_15_CLKBUF1_28 gnd vdd FILL
XFILL_24_DFFSR_125 gnd vdd FILL
XFILL_24_DFFSR_136 gnd vdd FILL
XFILL_15_CLKBUF1_39 gnd vdd FILL
XFILL_24_DFFSR_147 gnd vdd FILL
XFILL_10_AOI21X1_14 gnd vdd FILL
XFILL_24_DFFSR_158 gnd vdd FILL
XFILL_10_AOI21X1_25 gnd vdd FILL
XFILL_10_AOI21X1_36 gnd vdd FILL
XFILL_24_DFFSR_169 gnd vdd FILL
XFILL_10_AOI21X1_47 gnd vdd FILL
XFILL_1_DFFSR_13 gnd vdd FILL
XFILL_28_DFFSR_102 gnd vdd FILL
XFILL_5_INVX1_109 gnd vdd FILL
XFILL_1_DFFSR_24 gnd vdd FILL
XFILL_28_DFFSR_113 gnd vdd FILL
XFILL_10_AOI21X1_58 gnd vdd FILL
XFILL_1_DFFSR_35 gnd vdd FILL
XFILL_10_AOI21X1_69 gnd vdd FILL
XFILL_11_NOR2X1_1 gnd vdd FILL
XFILL_28_DFFSR_124 gnd vdd FILL
XFILL_28_DFFSR_135 gnd vdd FILL
XFILL_1_DFFSR_46 gnd vdd FILL
XFILL_28_DFFSR_146 gnd vdd FILL
XFILL_1_DFFSR_57 gnd vdd FILL
XFILL_28_DFFSR_157 gnd vdd FILL
XFILL_1_DFFSR_68 gnd vdd FILL
XFILL_1_DFFSR_79 gnd vdd FILL
XFILL_28_DFFSR_168 gnd vdd FILL
XFILL_28_DFFSR_179 gnd vdd FILL
XFILL_20_NOR3X1_15 gnd vdd FILL
XFILL_20_NOR3X1_26 gnd vdd FILL
XFILL_24_6_1 gnd vdd FILL
XFILL_20_NOR3X1_37 gnd vdd FILL
XFILL_20_NOR3X1_48 gnd vdd FILL
XFILL_70_DFFSR_204 gnd vdd FILL
XFILL_23_1_0 gnd vdd FILL
XFILL_70_DFFSR_215 gnd vdd FILL
XFILL_70_DFFSR_226 gnd vdd FILL
XFILL_12_NAND3X1_108 gnd vdd FILL
XFILL_70_DFFSR_237 gnd vdd FILL
XFILL_49_DFFSR_70 gnd vdd FILL
XFILL_70_DFFSR_248 gnd vdd FILL
XFILL_12_NAND3X1_119 gnd vdd FILL
XFILL_24_NOR3X1_14 gnd vdd FILL
XFILL_49_DFFSR_81 gnd vdd FILL
XFILL_70_DFFSR_259 gnd vdd FILL
XFILL_49_DFFSR_92 gnd vdd FILL
XFILL_24_NOR3X1_25 gnd vdd FILL
XFILL_24_NOR3X1_36 gnd vdd FILL
XFILL_24_NOR3X1_47 gnd vdd FILL
XFILL_74_DFFSR_203 gnd vdd FILL
XFILL_22_CLKBUF1_30 gnd vdd FILL
XFILL_74_DFFSR_214 gnd vdd FILL
XFILL_22_CLKBUF1_41 gnd vdd FILL
XFILL_74_DFFSR_225 gnd vdd FILL
XFILL_74_DFFSR_236 gnd vdd FILL
XFILL_74_DFFSR_247 gnd vdd FILL
XFILL_5_CLKBUF1_12 gnd vdd FILL
XFILL_28_NOR3X1_13 gnd vdd FILL
XFILL_74_DFFSR_258 gnd vdd FILL
XFILL_3_BUFX4_6 gnd vdd FILL
XFILL_74_DFFSR_269 gnd vdd FILL
XFILL_5_CLKBUF1_23 gnd vdd FILL
XFILL_28_NOR3X1_24 gnd vdd FILL
XFILL_5_CLKBUF1_34 gnd vdd FILL
XFILL_28_NOR3X1_35 gnd vdd FILL
XFILL_18_DFFSR_80 gnd vdd FILL
XFILL_78_DFFSR_202 gnd vdd FILL
XFILL_28_NOR3X1_46 gnd vdd FILL
XFILL_13_MUX2X1_108 gnd vdd FILL
XOAI22X1_6 INVX1_91/Y OAI22X1_6/B INVX1_94/Y OAI22X1_6/D gnd OAI22X1_6/Y vdd OAI22X1
XFILL_0_AOI21X1_20 gnd vdd FILL
XFILL_78_DFFSR_213 gnd vdd FILL
XFILL_13_MUX2X1_119 gnd vdd FILL
XFILL_18_DFFSR_91 gnd vdd FILL
XFILL_78_DFFSR_224 gnd vdd FILL
XFILL_78_DFFSR_235 gnd vdd FILL
XFILL_0_AOI21X1_31 gnd vdd FILL
XFILL_0_AOI21X1_42 gnd vdd FILL
XFILL_78_DFFSR_246 gnd vdd FILL
XFILL_0_AOI21X1_53 gnd vdd FILL
XFILL_10_OAI22X1_11 gnd vdd FILL
XFILL_0_AOI21X1_64 gnd vdd FILL
XFILL_78_DFFSR_257 gnd vdd FILL
XFILL_78_DFFSR_268 gnd vdd FILL
XFILL_0_AOI21X1_75 gnd vdd FILL
XFILL_10_OAI22X1_22 gnd vdd FILL
XFILL_33_CLKBUF1_9 gnd vdd FILL
XFILL_13_DFFSR_190 gnd vdd FILL
XFILL_10_OAI22X1_33 gnd vdd FILL
XFILL_10_OAI22X1_44 gnd vdd FILL
XFILL_58_DFFSR_90 gnd vdd FILL
XFILL_14_OAI21X1_13 gnd vdd FILL
XFILL_14_OAI21X1_24 gnd vdd FILL
XFILL_14_OAI21X1_35 gnd vdd FILL
XFILL_3_NOR2X1_130 gnd vdd FILL
XFILL_3_NOR2X1_141 gnd vdd FILL
XFILL_7_7_1 gnd vdd FILL
XFILL_14_OAI21X1_46 gnd vdd FILL
XFILL_3_NOR2X1_152 gnd vdd FILL
XFILL_6_2_0 gnd vdd FILL
XFILL_3_NOR2X1_163 gnd vdd FILL
XFILL_3_NOR2X1_174 gnd vdd FILL
XFILL_3_NOR2X1_185 gnd vdd FILL
XFILL_3_NOR2X1_196 gnd vdd FILL
XFILL_20_MUX2X1_110 gnd vdd FILL
XFILL_20_MUX2X1_121 gnd vdd FILL
XFILL_15_6_1 gnd vdd FILL
XFILL_20_MUX2X1_132 gnd vdd FILL
XFILL_20_MUX2X1_143 gnd vdd FILL
XFILL_20_MUX2X1_154 gnd vdd FILL
XFILL_14_1_0 gnd vdd FILL
XFILL_20_MUX2X1_165 gnd vdd FILL
XFILL_3_MUX2X1_103 gnd vdd FILL
XFILL_3_MUX2X1_114 gnd vdd FILL
XFILL_20_MUX2X1_176 gnd vdd FILL
XFILL_3_MUX2X1_125 gnd vdd FILL
XFILL_20_MUX2X1_187 gnd vdd FILL
XFILL_14_9 gnd vdd FILL
XFILL_3_MUX2X1_136 gnd vdd FILL
XFILL_14_BUFX4_18 gnd vdd FILL
XFILL_3_MUX2X1_147 gnd vdd FILL
XFILL_3_MUX2X1_158 gnd vdd FILL
XFILL_14_BUFX4_29 gnd vdd FILL
XFILL_3_MUX2X1_169 gnd vdd FILL
XFILL_6_INVX8_4 gnd vdd FILL
XDFFSR_208 INVX1_92/A CLKBUF1_7/Y BUFX4_13/Y vdd MUX2X1_78/Y gnd vdd DFFSR
XFILL_0_OAI22X1_50 gnd vdd FILL
XDFFSR_219 INVX1_77/A DFFSR_47/CLK DFFSR_6/R vdd MUX2X1_64/Y gnd vdd DFFSR
XFILL_19_INVX8_2 gnd vdd FILL
XFILL_4_OAI21X1_30 gnd vdd FILL
XFILL_41_DFFSR_203 gnd vdd FILL
XFILL_4_OAI21X1_41 gnd vdd FILL
XFILL_41_DFFSR_214 gnd vdd FILL
XFILL_3_OAI21X1_4 gnd vdd FILL
XFILL_41_DFFSR_225 gnd vdd FILL
XFILL_0_NOR2X1_40 gnd vdd FILL
XFILL_0_NOR2X1_51 gnd vdd FILL
XFILL_41_DFFSR_236 gnd vdd FILL
XFILL_0_NOR2X1_62 gnd vdd FILL
XFILL_41_DFFSR_247 gnd vdd FILL
XFILL_41_DFFSR_258 gnd vdd FILL
XFILL_41_DFFSR_269 gnd vdd FILL
XFILL_0_NOR2X1_73 gnd vdd FILL
XFILL_0_NOR2X1_84 gnd vdd FILL
XFILL_0_NOR2X1_95 gnd vdd FILL
XFILL_45_DFFSR_202 gnd vdd FILL
XFILL_23_DFFSR_4 gnd vdd FILL
XFILL_45_DFFSR_213 gnd vdd FILL
XFILL_7_OAI21X1_3 gnd vdd FILL
XFILL_45_DFFSR_224 gnd vdd FILL
XFILL_80_DFFSR_5 gnd vdd FILL
XFILL_45_DFFSR_235 gnd vdd FILL
XFILL_4_NOR2X1_50 gnd vdd FILL
XFILL_4_NOR2X1_61 gnd vdd FILL
XFILL_45_DFFSR_246 gnd vdd FILL
XFILL_45_DFFSR_257 gnd vdd FILL
XFILL_4_NOR2X1_72 gnd vdd FILL
XFILL_45_DFFSR_268 gnd vdd FILL
XFILL_4_NOR2X1_83 gnd vdd FILL
XFILL_72_DFFSR_102 gnd vdd FILL
XFILL_4_NOR2X1_94 gnd vdd FILL
XFILL_49_DFFSR_201 gnd vdd FILL
XFILL_49_DFFSR_212 gnd vdd FILL
XFILL_72_DFFSR_113 gnd vdd FILL
XFILL_72_DFFSR_124 gnd vdd FILL
XFILL_49_DFFSR_223 gnd vdd FILL
XFILL_49_DFFSR_234 gnd vdd FILL
XFILL_72_DFFSR_135 gnd vdd FILL
XFILL_72_DFFSR_146 gnd vdd FILL
XFILL_72_DFFSR_157 gnd vdd FILL
XFILL_8_NOR2X1_60 gnd vdd FILL
XFILL_49_DFFSR_245 gnd vdd FILL
XFILL_8_NOR2X1_71 gnd vdd FILL
XFILL_49_DFFSR_256 gnd vdd FILL
XFILL_49_DFFSR_267 gnd vdd FILL
XFILL_72_DFFSR_168 gnd vdd FILL
XFILL_65_5_1 gnd vdd FILL
XFILL_72_DFFSR_179 gnd vdd FILL
XFILL_8_NOR2X1_82 gnd vdd FILL
XFILL_76_DFFSR_101 gnd vdd FILL
XFILL_8_NOR2X1_93 gnd vdd FILL
XFILL_76_DFFSR_112 gnd vdd FILL
XFILL_64_0_0 gnd vdd FILL
XFILL_6_NAND3X1_17 gnd vdd FILL
XFILL_76_DFFSR_123 gnd vdd FILL
XFILL_76_DFFSR_134 gnd vdd FILL
XFILL_6_NAND3X1_28 gnd vdd FILL
XFILL_76_DFFSR_145 gnd vdd FILL
XFILL_6_NAND3X1_39 gnd vdd FILL
XFILL_76_DFFSR_156 gnd vdd FILL
XFILL_76_DFFSR_167 gnd vdd FILL
XFILL_76_DFFSR_178 gnd vdd FILL
XFILL_45_DFFSR_8 gnd vdd FILL
XFILL_6_BUFX4_17 gnd vdd FILL
XFILL_76_DFFSR_189 gnd vdd FILL
XFILL_6_BUFX4_28 gnd vdd FILL
XFILL_6_BUFX4_39 gnd vdd FILL
XFILL_0_NAND2X1_6 gnd vdd FILL
XFILL_4_NAND2X1_5 gnd vdd FILL
XFILL_0_MUX2X1_80 gnd vdd FILL
XFILL_13_AND2X2_5 gnd vdd FILL
XFILL_0_MUX2X1_91 gnd vdd FILL
XFILL_8_NAND2X1_4 gnd vdd FILL
XFILL_12_DFFSR_202 gnd vdd FILL
XFILL_12_DFFSR_213 gnd vdd FILL
XFILL_12_DFFSR_224 gnd vdd FILL
XFILL_12_DFFSR_235 gnd vdd FILL
XFILL_12_DFFSR_246 gnd vdd FILL
XFILL_4_MUX2X1_90 gnd vdd FILL
XFILL_12_DFFSR_257 gnd vdd FILL
XFILL_12_DFFSR_268 gnd vdd FILL
XFILL_10_BUFX4_11 gnd vdd FILL
XFILL_16_DFFSR_201 gnd vdd FILL
XFILL_25_CLKBUF1_18 gnd vdd FILL
XFILL_10_BUFX4_22 gnd vdd FILL
XFILL_16_DFFSR_212 gnd vdd FILL
XFILL_13_NAND3X1_1 gnd vdd FILL
XFILL_25_CLKBUF1_29 gnd vdd FILL
XFILL_10_BUFX4_33 gnd vdd FILL
XFILL_16_DFFSR_223 gnd vdd FILL
XFILL_10_BUFX4_44 gnd vdd FILL
XFILL_56_5_1 gnd vdd FILL
XFILL_16_DFFSR_234 gnd vdd FILL
XFILL_10_BUFX4_55 gnd vdd FILL
XFILL_16_DFFSR_245 gnd vdd FILL
XFILL_55_0_0 gnd vdd FILL
XFILL_16_DFFSR_256 gnd vdd FILL
XFILL_10_BUFX4_66 gnd vdd FILL
XFILL_7_BUFX4_7 gnd vdd FILL
XFILL_16_DFFSR_267 gnd vdd FILL
XFILL_10_BUFX4_77 gnd vdd FILL
XFILL_10_BUFX4_88 gnd vdd FILL
XFILL_43_DFFSR_101 gnd vdd FILL
XFILL_10_BUFX4_99 gnd vdd FILL
XFILL_43_DFFSR_112 gnd vdd FILL
XFILL_3_AOI21X1_19 gnd vdd FILL
XFILL_43_DFFSR_123 gnd vdd FILL
XFILL_43_DFFSR_134 gnd vdd FILL
XFILL_43_DFFSR_145 gnd vdd FILL
XFILL_43_DFFSR_156 gnd vdd FILL
XFILL_43_DFFSR_167 gnd vdd FILL
XFILL_43_DFFSR_178 gnd vdd FILL
XFILL_47_DFFSR_100 gnd vdd FILL
XFILL_43_DFFSR_189 gnd vdd FILL
XFILL_47_DFFSR_111 gnd vdd FILL
XFILL_6_NOR2X1_107 gnd vdd FILL
XFILL_47_DFFSR_122 gnd vdd FILL
XFILL_6_NOR2X1_118 gnd vdd FILL
XFILL_8_AOI21X1_9 gnd vdd FILL
XFILL_47_DFFSR_133 gnd vdd FILL
XFILL_47_DFFSR_144 gnd vdd FILL
XFILL_6_NOR2X1_129 gnd vdd FILL
XFILL_12_NAND3X1_20 gnd vdd FILL
XFILL_47_DFFSR_155 gnd vdd FILL
XFILL_12_NAND3X1_31 gnd vdd FILL
XFILL_47_DFFSR_166 gnd vdd FILL
XFILL_13_NAND3X1_109 gnd vdd FILL
XFILL_47_DFFSR_177 gnd vdd FILL
XFILL_12_NAND3X1_42 gnd vdd FILL
XFILL_4_INVX1_12 gnd vdd FILL
XFILL_12_NAND3X1_53 gnd vdd FILL
XFILL_4_INVX1_23 gnd vdd FILL
XFILL_47_DFFSR_188 gnd vdd FILL
XFILL_4_INVX1_34 gnd vdd FILL
XFILL_12_NAND3X1_64 gnd vdd FILL
XFILL_47_DFFSR_199 gnd vdd FILL
XFILL_32_CLKBUF1_20 gnd vdd FILL
XFILL_12_NAND3X1_75 gnd vdd FILL
XFILL_5_AND2X2_4 gnd vdd FILL
XFILL_12_NAND3X1_86 gnd vdd FILL
XFILL_4_INVX1_45 gnd vdd FILL
XFILL_4_INVX1_56 gnd vdd FILL
XFILL_32_CLKBUF1_31 gnd vdd FILL
XFILL_12_NAND3X1_97 gnd vdd FILL
XFILL_4_INVX1_67 gnd vdd FILL
XFILL_32_CLKBUF1_42 gnd vdd FILL
XFILL_3_BUFX2_3 gnd vdd FILL
XFILL_13_AOI22X1_6 gnd vdd FILL
XFILL_4_INVX1_78 gnd vdd FILL
XFILL_4_INVX1_89 gnd vdd FILL
XFILL_23_MUX2X1_109 gnd vdd FILL
XFILL_17_AOI22X1_5 gnd vdd FILL
XFILL_2_BUFX4_10 gnd vdd FILL
XFILL_2_BUFX4_21 gnd vdd FILL
XFILL_62_DFFSR_2 gnd vdd FILL
XFILL_2_BUFX4_32 gnd vdd FILL
XFILL_2_BUFX4_43 gnd vdd FILL
XFILL_19_DFFSR_14 gnd vdd FILL
XFILL_2_BUFX4_54 gnd vdd FILL
XFILL_2_BUFX4_65 gnd vdd FILL
XFILL_19_DFFSR_25 gnd vdd FILL
XFILL_2_BUFX4_76 gnd vdd FILL
XFILL_19_DFFSR_36 gnd vdd FILL
XFILL_19_DFFSR_47 gnd vdd FILL
XFILL_19_DFFSR_58 gnd vdd FILL
XFILL_2_BUFX4_87 gnd vdd FILL
XFILL_3_OAI22X1_16 gnd vdd FILL
XFILL_19_DFFSR_69 gnd vdd FILL
XFILL_3_OAI22X1_27 gnd vdd FILL
XFILL_2_BUFX4_98 gnd vdd FILL
XFILL_3_OAI22X1_38 gnd vdd FILL
XFILL_3_OAI22X1_49 gnd vdd FILL
XFILL_59_DFFSR_13 gnd vdd FILL
XFILL_47_5_1 gnd vdd FILL
XFILL_59_DFFSR_24 gnd vdd FILL
XFILL_7_OAI21X1_18 gnd vdd FILL
XFILL_7_OAI21X1_29 gnd vdd FILL
XFILL_59_DFFSR_35 gnd vdd FILL
XFILL_46_0_0 gnd vdd FILL
XFILL_59_DFFSR_46 gnd vdd FILL
XFILL_59_DFFSR_57 gnd vdd FILL
XFILL_59_DFFSR_68 gnd vdd FILL
XFILL_20_MUX2X1_8 gnd vdd FILL
XFILL_59_DFFSR_79 gnd vdd FILL
XFILL_2_NAND3X1_70 gnd vdd FILL
XFILL_10_DFFSR_101 gnd vdd FILL
XFILL_2_NAND3X1_81 gnd vdd FILL
XFILL_2_NAND3X1_92 gnd vdd FILL
XFILL_27_DFFSR_5 gnd vdd FILL
XFILL_6_NAND2X1_50 gnd vdd FILL
XFILL_10_DFFSR_112 gnd vdd FILL
XFILL_6_NAND2X1_61 gnd vdd FILL
XFILL_10_DFFSR_123 gnd vdd FILL
XFILL_10_DFFSR_134 gnd vdd FILL
XFILL_84_DFFSR_6 gnd vdd FILL
XFILL_6_NAND2X1_72 gnd vdd FILL
XFILL_28_DFFSR_12 gnd vdd FILL
XFILL_10_DFFSR_145 gnd vdd FILL
XFILL_6_NAND2X1_83 gnd vdd FILL
XFILL_10_DFFSR_156 gnd vdd FILL
XFILL_28_DFFSR_23 gnd vdd FILL
XFILL_6_NAND2X1_94 gnd vdd FILL
XFILL_28_DFFSR_34 gnd vdd FILL
XFILL_10_DFFSR_167 gnd vdd FILL
XFILL_3_INVX2_3 gnd vdd FILL
XFILL_10_DFFSR_178 gnd vdd FILL
XFILL_28_DFFSR_45 gnd vdd FILL
XFILL_28_DFFSR_56 gnd vdd FILL
XFILL_14_DFFSR_100 gnd vdd FILL
XFILL_10_DFFSR_189 gnd vdd FILL
XFILL_30_4_1 gnd vdd FILL
XFILL_28_DFFSR_67 gnd vdd FILL
XFILL_14_DFFSR_111 gnd vdd FILL
XFILL_14_CLKBUF1_14 gnd vdd FILL
XFILL_28_DFFSR_78 gnd vdd FILL
XFILL_28_DFFSR_89 gnd vdd FILL
XFILL_14_CLKBUF1_25 gnd vdd FILL
XFILL_14_DFFSR_122 gnd vdd FILL
XFILL_14_CLKBUF1_36 gnd vdd FILL
XFILL_14_DFFSR_133 gnd vdd FILL
XFILL_14_DFFSR_144 gnd vdd FILL
XFILL_68_DFFSR_11 gnd vdd FILL
XFILL_14_DFFSR_155 gnd vdd FILL
XFILL_68_DFFSR_22 gnd vdd FILL
XFILL_68_DFFSR_33 gnd vdd FILL
XFILL_14_DFFSR_166 gnd vdd FILL
XFILL_68_DFFSR_44 gnd vdd FILL
XFILL_3_CLKBUF1_9 gnd vdd FILL
XFILL_14_DFFSR_177 gnd vdd FILL
XFILL_3_MUX2X1_9 gnd vdd FILL
XFILL_68_DFFSR_55 gnd vdd FILL
XFILL_14_DFFSR_188 gnd vdd FILL
XFILL_68_DFFSR_66 gnd vdd FILL
XFILL_18_DFFSR_110 gnd vdd FILL
XFILL_14_DFFSR_199 gnd vdd FILL
XFILL_68_DFFSR_77 gnd vdd FILL
XFILL_1_INVX1_1 gnd vdd FILL
XFILL_68_DFFSR_88 gnd vdd FILL
XFILL_18_DFFSR_121 gnd vdd FILL
XFILL_18_DFFSR_132 gnd vdd FILL
XFILL_68_DFFSR_99 gnd vdd FILL
XFILL_18_DFFSR_143 gnd vdd FILL
XFILL_18_DFFSR_154 gnd vdd FILL
XFILL_18_DFFSR_165 gnd vdd FILL
XFILL_49_DFFSR_9 gnd vdd FILL
XFILL_7_CLKBUF1_8 gnd vdd FILL
XFILL_10_NOR3X1_12 gnd vdd FILL
XFILL_18_DFFSR_176 gnd vdd FILL
XFILL_18_DFFSR_187 gnd vdd FILL
XFILL_10_NOR3X1_23 gnd vdd FILL
XFILL_37_DFFSR_10 gnd vdd FILL
XFILL_10_NOR3X1_34 gnd vdd FILL
XFILL_37_DFFSR_21 gnd vdd FILL
XFILL_18_DFFSR_198 gnd vdd FILL
XFILL_37_DFFSR_32 gnd vdd FILL
XFILL_60_DFFSR_201 gnd vdd FILL
XFILL_37_DFFSR_43 gnd vdd FILL
XFILL_10_NOR3X1_45 gnd vdd FILL
XFILL_60_DFFSR_212 gnd vdd FILL
XFILL_37_DFFSR_54 gnd vdd FILL
XFILL_60_DFFSR_223 gnd vdd FILL
XFILL_37_DFFSR_65 gnd vdd FILL
XFILL_3_BUFX4_103 gnd vdd FILL
XFILL_37_DFFSR_76 gnd vdd FILL
XFILL_60_DFFSR_234 gnd vdd FILL
XFILL_37_DFFSR_87 gnd vdd FILL
XFILL_60_DFFSR_245 gnd vdd FILL
XFILL_14_NOR3X1_11 gnd vdd FILL
XFILL_37_DFFSR_98 gnd vdd FILL
XFILL_60_DFFSR_256 gnd vdd FILL
XFILL_60_DFFSR_267 gnd vdd FILL
XFILL_14_NOR3X1_22 gnd vdd FILL
XFILL_14_NOR3X1_33 gnd vdd FILL
XFILL_77_DFFSR_20 gnd vdd FILL
XFILL_77_DFFSR_31 gnd vdd FILL
XFILL_64_DFFSR_200 gnd vdd FILL
XFILL_14_NOR3X1_44 gnd vdd FILL
XFILL_77_DFFSR_42 gnd vdd FILL
XFILL_64_DFFSR_211 gnd vdd FILL
XFILL_77_DFFSR_53 gnd vdd FILL
XFILL_64_DFFSR_222 gnd vdd FILL
XFILL_77_DFFSR_64 gnd vdd FILL
XFILL_64_DFFSR_233 gnd vdd FILL
XFILL_7_BUFX4_102 gnd vdd FILL
XFILL_38_5_1 gnd vdd FILL
XFILL_77_DFFSR_75 gnd vdd FILL
XFILL_77_DFFSR_86 gnd vdd FILL
XFILL_64_DFFSR_244 gnd vdd FILL
XFILL_18_NOR3X1_10 gnd vdd FILL
XFILL_37_0_0 gnd vdd FILL
XFILL_64_DFFSR_255 gnd vdd FILL
XFILL_77_DFFSR_97 gnd vdd FILL
XFILL_4_CLKBUF1_20 gnd vdd FILL
XFILL_64_DFFSR_266 gnd vdd FILL
XFILL_18_NOR3X1_21 gnd vdd FILL
XFILL_4_CLKBUF1_31 gnd vdd FILL
XFILL_18_NOR3X1_32 gnd vdd FILL
XFILL_4_CLKBUF1_42 gnd vdd FILL
XFILL_18_NOR3X1_43 gnd vdd FILL
XFILL_0_INVX1_60 gnd vdd FILL
XFILL_12_MUX2X1_105 gnd vdd FILL
XFILL_68_DFFSR_210 gnd vdd FILL
XFILL_0_INVX1_71 gnd vdd FILL
XFILL_0_INVX1_82 gnd vdd FILL
XFILL_12_MUX2X1_116 gnd vdd FILL
XFILL_68_DFFSR_221 gnd vdd FILL
XFILL_0_INVX1_93 gnd vdd FILL
XFILL_12_MUX2X1_127 gnd vdd FILL
XFILL_68_DFFSR_232 gnd vdd FILL
XFILL_12_MUX2X1_138 gnd vdd FILL
XFILL_46_DFFSR_30 gnd vdd FILL
XFILL_68_DFFSR_243 gnd vdd FILL
XFILL_12_MUX2X1_149 gnd vdd FILL
XFILL_46_DFFSR_41 gnd vdd FILL
XFILL_17_NOR3X1_5 gnd vdd FILL
XFILL_68_DFFSR_254 gnd vdd FILL
XFILL_46_DFFSR_52 gnd vdd FILL
XFILL_46_DFFSR_63 gnd vdd FILL
XFILL_68_DFFSR_265 gnd vdd FILL
XFILL_46_DFFSR_74 gnd vdd FILL
XFILL_23_CLKBUF1_6 gnd vdd FILL
XFILL_46_DFFSR_85 gnd vdd FILL
XFILL_13_OAI21X1_10 gnd vdd FILL
XFILL_46_DFFSR_96 gnd vdd FILL
XFILL_1_NOR2X1_16 gnd vdd FILL
XFILL_13_OAI21X1_21 gnd vdd FILL
XFILL_1_NOR2X1_27 gnd vdd FILL
XFILL_13_OAI21X1_32 gnd vdd FILL
XFILL_1_NOR2X1_38 gnd vdd FILL
XFILL_13_OAI21X1_43 gnd vdd FILL
XFILL_21_4_1 gnd vdd FILL
XFILL_1_NOR2X1_49 gnd vdd FILL
XFILL_86_DFFSR_40 gnd vdd FILL
XFILL_2_NOR2X1_160 gnd vdd FILL
XFILL_86_DFFSR_51 gnd vdd FILL
XFILL_86_DFFSR_62 gnd vdd FILL
XFILL_2_NOR2X1_171 gnd vdd FILL
XFILL_86_DFFSR_73 gnd vdd FILL
XFILL_27_CLKBUF1_5 gnd vdd FILL
XFILL_86_DFFSR_84 gnd vdd FILL
XFILL_2_NOR2X1_182 gnd vdd FILL
XFILL_15_DFFSR_40 gnd vdd FILL
XFILL_2_NOR2X1_193 gnd vdd FILL
XFILL_5_NOR2X1_15 gnd vdd FILL
XFILL_86_DFFSR_95 gnd vdd FILL
XFILL_15_DFFSR_51 gnd vdd FILL
XFILL_5_NOR2X1_26 gnd vdd FILL
XFILL_15_DFFSR_62 gnd vdd FILL
XFILL_5_NOR2X1_37 gnd vdd FILL
XFILL_15_DFFSR_73 gnd vdd FILL
XFILL_15_DFFSR_84 gnd vdd FILL
XFILL_5_NOR2X1_48 gnd vdd FILL
XFILL_5_NOR2X1_59 gnd vdd FILL
XFILL_15_DFFSR_95 gnd vdd FILL
XFILL_26_NOR3X1_3 gnd vdd FILL
XFILL_9_NOR2X1_14 gnd vdd FILL
XFILL_9_NOR2X1_25 gnd vdd FILL
XFILL_55_DFFSR_50 gnd vdd FILL
XFILL_55_DFFSR_61 gnd vdd FILL
XFILL_9_NOR2X1_36 gnd vdd FILL
XFILL_55_DFFSR_72 gnd vdd FILL
XFILL_55_DFFSR_83 gnd vdd FILL
XFILL_9_NOR2X1_47 gnd vdd FILL
XFILL_9_NOR2X1_58 gnd vdd FILL
XFILL_55_DFFSR_94 gnd vdd FILL
XFILL_13_OAI22X1_9 gnd vdd FILL
XFILL_9_NOR2X1_69 gnd vdd FILL
XFILL_2_MUX2X1_100 gnd vdd FILL
XFILL_2_MUX2X1_111 gnd vdd FILL
XFILL_0_NOR2X1_4 gnd vdd FILL
XFILL_2_MUX2X1_122 gnd vdd FILL
XFILL_2_MUX2X1_133 gnd vdd FILL
XFILL_2_MUX2X1_144 gnd vdd FILL
XFILL_2_MUX2X1_155 gnd vdd FILL
XFILL_15_NAND3X1_19 gnd vdd FILL
XFILL_17_OAI22X1_8 gnd vdd FILL
XFILL_2_MUX2X1_166 gnd vdd FILL
XFILL_2_MUX2X1_177 gnd vdd FILL
XFILL_2_MUX2X1_188 gnd vdd FILL
XFILL_24_DFFSR_60 gnd vdd FILL
XFILL_24_DFFSR_71 gnd vdd FILL
XFILL_24_DFFSR_82 gnd vdd FILL
XFILL_24_DFFSR_93 gnd vdd FILL
XFILL_4_5_1 gnd vdd FILL
XFILL_29_5_1 gnd vdd FILL
XFILL_35_CLKBUF1_19 gnd vdd FILL
XFILL_31_DFFSR_200 gnd vdd FILL
XFILL_9_NOR3X1_4 gnd vdd FILL
XFILL_31_DFFSR_211 gnd vdd FILL
XFILL_28_0_0 gnd vdd FILL
XFILL_31_DFFSR_222 gnd vdd FILL
XFILL_3_0_0 gnd vdd FILL
XFILL_7_BUFX2_4 gnd vdd FILL
XFILL_31_DFFSR_233 gnd vdd FILL
XFILL_31_DFFSR_244 gnd vdd FILL
XFILL_31_DFFSR_255 gnd vdd FILL
XFILL_64_DFFSR_70 gnd vdd FILL
XFILL_31_DFFSR_266 gnd vdd FILL
XFILL_64_DFFSR_81 gnd vdd FILL
XFILL_64_DFFSR_92 gnd vdd FILL
XFILL_35_DFFSR_210 gnd vdd FILL
XFILL_35_DFFSR_221 gnd vdd FILL
XFILL_35_DFFSR_232 gnd vdd FILL
XFILL_35_DFFSR_243 gnd vdd FILL
XFILL_66_DFFSR_3 gnd vdd FILL
XFILL_35_DFFSR_254 gnd vdd FILL
XFILL_7_DFFSR_50 gnd vdd FILL
XFILL_1_MUX2X1_12 gnd vdd FILL
XFILL_35_DFFSR_265 gnd vdd FILL
XFILL_7_DFFSR_61 gnd vdd FILL
XFILL_1_MUX2X1_23 gnd vdd FILL
XFILL_12_4_1 gnd vdd FILL
XFILL_7_DFFSR_72 gnd vdd FILL
XFILL_7_DFFSR_83 gnd vdd FILL
XFILL_1_MUX2X1_34 gnd vdd FILL
XFILL_62_DFFSR_110 gnd vdd FILL
XINVX8_2 din[2] gnd INVX8_2/Y vdd INVX8
XFILL_1_MUX2X1_45 gnd vdd FILL
XFILL_7_DFFSR_94 gnd vdd FILL
XFILL_39_DFFSR_220 gnd vdd FILL
XFILL_62_DFFSR_121 gnd vdd FILL
XFILL_1_MUX2X1_56 gnd vdd FILL
XFILL_33_DFFSR_80 gnd vdd FILL
XFILL_62_DFFSR_132 gnd vdd FILL
XFILL_39_DFFSR_231 gnd vdd FILL
XFILL_1_MUX2X1_67 gnd vdd FILL
XFILL_62_DFFSR_143 gnd vdd FILL
XFILL_39_DFFSR_242 gnd vdd FILL
XFILL_33_DFFSR_91 gnd vdd FILL
XFILL_62_DFFSR_154 gnd vdd FILL
XFILL_1_MUX2X1_78 gnd vdd FILL
XFILL_62_DFFSR_165 gnd vdd FILL
XFILL_39_DFFSR_253 gnd vdd FILL
XFILL_1_MUX2X1_89 gnd vdd FILL
XFILL_39_DFFSR_264 gnd vdd FILL
XFILL_5_MUX2X1_11 gnd vdd FILL
XFILL_39_DFFSR_275 gnd vdd FILL
XFILL_5_MUX2X1_22 gnd vdd FILL
XFILL_62_DFFSR_176 gnd vdd FILL
XFILL_62_DFFSR_187 gnd vdd FILL
XFILL_62_DFFSR_198 gnd vdd FILL
XFILL_5_MUX2X1_33 gnd vdd FILL
XFILL_66_DFFSR_120 gnd vdd FILL
XFILL_5_MUX2X1_44 gnd vdd FILL
XFILL_5_NAND3X1_14 gnd vdd FILL
XFILL_5_MUX2X1_55 gnd vdd FILL
XFILL_66_DFFSR_131 gnd vdd FILL
XFILL_5_NAND3X1_25 gnd vdd FILL
XFILL_5_MUX2X1_66 gnd vdd FILL
XFILL_73_DFFSR_90 gnd vdd FILL
XFILL_66_DFFSR_142 gnd vdd FILL
XFILL_5_NAND3X1_36 gnd vdd FILL
XFILL_5_MUX2X1_77 gnd vdd FILL
XFILL_66_DFFSR_153 gnd vdd FILL
XFILL_5_NAND3X1_47 gnd vdd FILL
XFILL_5_MUX2X1_88 gnd vdd FILL
XFILL_5_NAND3X1_58 gnd vdd FILL
XFILL_66_DFFSR_164 gnd vdd FILL
XFILL_5_MUX2X1_99 gnd vdd FILL
XFILL_50_DFFSR_9 gnd vdd FILL
XFILL_9_MUX2X1_10 gnd vdd FILL
XFILL_9_NAND2X1_16 gnd vdd FILL
XFILL_9_MUX2X1_21 gnd vdd FILL
XFILL_5_NAND3X1_69 gnd vdd FILL
XFILL_66_DFFSR_175 gnd vdd FILL
XFILL_9_NAND2X1_27 gnd vdd FILL
XFILL_66_DFFSR_186 gnd vdd FILL
XFILL_9_MUX2X1_32 gnd vdd FILL
XFILL_9_NAND2X1_38 gnd vdd FILL
XFILL_66_DFFSR_197 gnd vdd FILL
XFILL_9_NAND2X1_49 gnd vdd FILL
XFILL_9_MUX2X1_43 gnd vdd FILL
XFILL_9_MUX2X1_54 gnd vdd FILL
XFILL_9_MUX2X1_65 gnd vdd FILL
XFILL_9_MUX2X1_76 gnd vdd FILL
XFILL_9_MUX2X1_87 gnd vdd FILL
XFILL_9_MUX2X1_98 gnd vdd FILL
XFILL_7_INVX2_4 gnd vdd FILL
XBUFX4_11 BUFX4_44/A gnd DFFSR_90/R vdd BUFX4
XBUFX4_22 BUFX4_54/A gnd DFFSR_6/R vdd BUFX4
XFILL_19_MUX2X1_180 gnd vdd FILL
XBUFX4_33 BUFX4_47/A gnd DFFSR_4/R vdd BUFX4
XFILL_19_MUX2X1_191 gnd vdd FILL
XBUFX4_44 BUFX4_44/A gnd DFFSR_42/R vdd BUFX4
XBUFX4_55 BUFX4_62/Y gnd BUFX4_55/Y vdd BUFX4
XBUFX4_66 INVX8_1/Y gnd BUFX4_66/Y vdd BUFX4
XBUFX4_77 INVX8_2/Y gnd BUFX4_77/Y vdd BUFX4
XFILL_19_0_0 gnd vdd FILL
XBUFX4_88 BUFX4_92/A gnd BUFX4_88/Y vdd BUFX4
XBUFX4_99 INVX8_3/Y gnd BUFX4_99/Y vdd BUFX4
XFILL_48_DFFSR_109 gnd vdd FILL
XFILL_5_INVX1_2 gnd vdd FILL
XFILL_21_MUX2X1_20 gnd vdd FILL
XFILL_21_MUX2X1_31 gnd vdd FILL
XFILL_21_MUX2X1_42 gnd vdd FILL
XFILL_21_MUX2X1_53 gnd vdd FILL
XFILL_62_3_1 gnd vdd FILL
XFILL_21_MUX2X1_64 gnd vdd FILL
XFILL_21_MUX2X1_75 gnd vdd FILL
XFILL_21_MUX2X1_86 gnd vdd FILL
XFILL_21_MUX2X1_97 gnd vdd FILL
XFILL_10_3 gnd vdd FILL
XFILL_24_CLKBUF1_15 gnd vdd FILL
XFILL_24_CLKBUF1_26 gnd vdd FILL
XFILL_24_CLKBUF1_37 gnd vdd FILL
XFILL_7_CLKBUF1_19 gnd vdd FILL
XFILL_2_AOI21X1_16 gnd vdd FILL
XFILL_33_DFFSR_120 gnd vdd FILL
XFILL_33_DFFSR_131 gnd vdd FILL
XFILL_2_AOI21X1_27 gnd vdd FILL
XFILL_33_DFFSR_142 gnd vdd FILL
XFILL_33_DFFSR_153 gnd vdd FILL
XFILL_2_AOI21X1_38 gnd vdd FILL
XFILL_2_AOI21X1_49 gnd vdd FILL
XFILL_33_DFFSR_164 gnd vdd FILL
XFILL_33_DFFSR_175 gnd vdd FILL
XFILL_12_OAI22X1_18 gnd vdd FILL
XFILL_33_DFFSR_186 gnd vdd FILL
XFILL_12_OAI22X1_29 gnd vdd FILL
XFILL_33_DFFSR_197 gnd vdd FILL
XFILL_5_NOR2X1_104 gnd vdd FILL
XFILL_5_NOR2X1_115 gnd vdd FILL
XFILL_37_DFFSR_130 gnd vdd FILL
XFILL_5_NOR2X1_126 gnd vdd FILL
XFILL_37_DFFSR_141 gnd vdd FILL
XFILL_37_DFFSR_152 gnd vdd FILL
XFILL_5_NOR2X1_137 gnd vdd FILL
XFILL_37_DFFSR_163 gnd vdd FILL
XFILL_5_NOR2X1_148 gnd vdd FILL
XFILL_5_NOR2X1_159 gnd vdd FILL
XFILL_37_DFFSR_174 gnd vdd FILL
XFILL_11_NAND3X1_50 gnd vdd FILL
XFILL_37_DFFSR_185 gnd vdd FILL
XFILL_11_NAND3X1_61 gnd vdd FILL
XFILL_37_DFFSR_196 gnd vdd FILL
XFILL_11_NAND3X1_72 gnd vdd FILL
XFILL_11_NAND3X1_83 gnd vdd FILL
XFILL_11_NAND3X1_94 gnd vdd FILL
XFILL_15_DFFSR_109 gnd vdd FILL
XFILL_53_3_1 gnd vdd FILL
XFILL_22_MUX2X1_106 gnd vdd FILL
XFILL_22_MUX2X1_117 gnd vdd FILL
XFILL_83_DFFSR_220 gnd vdd FILL
XFILL_10_AOI21X1_5 gnd vdd FILL
XFILL_10_DFFSR_2 gnd vdd FILL
XFILL_22_MUX2X1_128 gnd vdd FILL
XFILL_83_DFFSR_231 gnd vdd FILL
XFILL_22_MUX2X1_139 gnd vdd FILL
XFILL_83_DFFSR_242 gnd vdd FILL
XFILL_83_DFFSR_253 gnd vdd FILL
XFILL_83_DFFSR_264 gnd vdd FILL
XFILL_83_DFFSR_275 gnd vdd FILL
XFILL_19_DFFSR_108 gnd vdd FILL
XFILL_19_DFFSR_119 gnd vdd FILL
XFILL_1_INVX1_16 gnd vdd FILL
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XFILL_1_INVX1_27 gnd vdd FILL
XFILL_1_INVX1_38 gnd vdd FILL
XFILL_87_DFFSR_230 gnd vdd FILL
XFILL_14_AOI21X1_4 gnd vdd FILL
XFILL_2_OAI22X1_13 gnd vdd FILL
XFILL_87_DFFSR_241 gnd vdd FILL
XFILL_2_AND2X2_8 gnd vdd FILL
XFILL_1_INVX1_49 gnd vdd FILL
XFILL_2_OAI22X1_24 gnd vdd FILL
XFILL_2_OAI22X1_35 gnd vdd FILL
XFILL_87_DFFSR_252 gnd vdd FILL
XFILL_2_OAI22X1_46 gnd vdd FILL
XFILL_87_DFFSR_263 gnd vdd FILL
XFILL_87_DFFSR_274 gnd vdd FILL
XFILL_47_DFFSR_19 gnd vdd FILL
XFILL_6_OAI21X1_15 gnd vdd FILL
XFILL_6_OAI21X1_26 gnd vdd FILL
XFILL_6_OAI21X1_37 gnd vdd FILL
XFILL_6_OAI21X1_48 gnd vdd FILL
XFILL_3_INVX1_180 gnd vdd FILL
XFILL_87_DFFSR_18 gnd vdd FILL
XFILL_3_INVX1_191 gnd vdd FILL
XFILL_32_DFFSR_6 gnd vdd FILL
XFILL_87_DFFSR_29 gnd vdd FILL
XFILL_65_DFFSR_209 gnd vdd FILL
XFILL_16_DFFSR_18 gnd vdd FILL
XFILL_5_NAND2X1_80 gnd vdd FILL
XFILL_5_NAND2X1_91 gnd vdd FILL
XFILL_16_DFFSR_29 gnd vdd FILL
XFILL_7_INVX1_190 gnd vdd FILL
XFILL_19_NOR3X1_19 gnd vdd FILL
XFILL_13_CLKBUF1_11 gnd vdd FILL
XFILL_9_OR2X2_1 gnd vdd FILL
XFILL_13_CLKBUF1_22 gnd vdd FILL
XFILL_69_DFFSR_208 gnd vdd FILL
XFILL_69_DFFSR_219 gnd vdd FILL
XFILL_13_CLKBUF1_33 gnd vdd FILL
XFILL_56_DFFSR_17 gnd vdd FILL
XFILL_56_DFFSR_28 gnd vdd FILL
XFILL_56_DFFSR_39 gnd vdd FILL
XFILL_44_3_1 gnd vdd FILL
XFILL_25_DFFSR_16 gnd vdd FILL
XFILL_11_NOR2X1_140 gnd vdd FILL
XFILL_11_NOR2X1_151 gnd vdd FILL
XFILL_25_DFFSR_27 gnd vdd FILL
XFILL_25_DFFSR_38 gnd vdd FILL
XFILL_11_NOR2X1_162 gnd vdd FILL
XFILL_11_NOR2X1_173 gnd vdd FILL
XFILL_25_DFFSR_49 gnd vdd FILL
XFILL_11_NOR2X1_184 gnd vdd FILL
XFILL_50_DFFSR_220 gnd vdd FILL
XFILL_11_NOR2X1_195 gnd vdd FILL
XFILL_50_DFFSR_231 gnd vdd FILL
XFILL_50_DFFSR_242 gnd vdd FILL
XFILL_50_DFFSR_253 gnd vdd FILL
XFILL_65_DFFSR_15 gnd vdd FILL
XFILL_65_DFFSR_26 gnd vdd FILL
XFILL_50_DFFSR_264 gnd vdd FILL
XFILL_50_DFFSR_275 gnd vdd FILL
XFILL_65_DFFSR_37 gnd vdd FILL
XFILL_65_DFFSR_48 gnd vdd FILL
XFILL_9_AOI21X1_80 gnd vdd FILL
XFILL_65_DFFSR_59 gnd vdd FILL
XFILL_54_DFFSR_230 gnd vdd FILL
XFILL_54_DFFSR_241 gnd vdd FILL
XFILL_54_DFFSR_252 gnd vdd FILL
XFILL_54_DFFSR_263 gnd vdd FILL
XFILL_54_DFFSR_274 gnd vdd FILL
XFILL_8_DFFSR_17 gnd vdd FILL
XFILL_8_DFFSR_28 gnd vdd FILL
XFILL_11_MUX2X1_102 gnd vdd FILL
XFILL_8_DFFSR_39 gnd vdd FILL
XFILL_11_MUX2X1_113 gnd vdd FILL
XFILL_34_DFFSR_14 gnd vdd FILL
XFILL_34_DFFSR_25 gnd vdd FILL
XFILL_81_DFFSR_130 gnd vdd FILL
XFILL_11_MUX2X1_124 gnd vdd FILL
XFILL_34_DFFSR_36 gnd vdd FILL
XFILL_11_MUX2X1_135 gnd vdd FILL
XFILL_58_DFFSR_240 gnd vdd FILL
XFILL_81_DFFSR_141 gnd vdd FILL
XFILL_34_DFFSR_47 gnd vdd FILL
XFILL_81_DFFSR_152 gnd vdd FILL
XFILL_11_MUX2X1_146 gnd vdd FILL
XFILL_34_DFFSR_58 gnd vdd FILL
XFILL_58_DFFSR_251 gnd vdd FILL
XFILL_81_DFFSR_163 gnd vdd FILL
XFILL_11_MUX2X1_157 gnd vdd FILL
XFILL_58_DFFSR_262 gnd vdd FILL
XFILL_34_DFFSR_69 gnd vdd FILL
XFILL_11_MUX2X1_168 gnd vdd FILL
XFILL_81_DFFSR_174 gnd vdd FILL
XFILL_13_CLKBUF1_3 gnd vdd FILL
XFILL_58_DFFSR_273 gnd vdd FILL
XFILL_1_DFFSR_200 gnd vdd FILL
XFILL_81_DFFSR_185 gnd vdd FILL
XFILL_11_MUX2X1_179 gnd vdd FILL
XFILL_74_DFFSR_13 gnd vdd FILL
XFILL_1_DFFSR_211 gnd vdd FILL
XFILL_81_DFFSR_196 gnd vdd FILL
XFILL_1_DFFSR_222 gnd vdd FILL
XFILL_32_DFFSR_209 gnd vdd FILL
XFILL_1_DFFSR_233 gnd vdd FILL
XFILL_74_DFFSR_24 gnd vdd FILL
XFILL_74_DFFSR_35 gnd vdd FILL
XFILL_9_2 gnd vdd FILL
XFILL_85_DFFSR_140 gnd vdd FILL
XFILL_74_DFFSR_46 gnd vdd FILL
XFILL_1_DFFSR_244 gnd vdd FILL
XFILL_12_OAI21X1_40 gnd vdd FILL
XFILL_74_DFFSR_57 gnd vdd FILL
XFILL_85_DFFSR_151 gnd vdd FILL
XFILL_1_DFFSR_255 gnd vdd FILL
XFILL_17_MUX2X1_3 gnd vdd FILL
XFILL_85_DFFSR_162 gnd vdd FILL
XFILL_74_DFFSR_68 gnd vdd FILL
XFILL_1_DFFSR_266 gnd vdd FILL
XFILL_85_DFFSR_173 gnd vdd FILL
XFILL_65_4 gnd vdd FILL
XFILL_74_DFFSR_79 gnd vdd FILL
XFILL_17_CLKBUF1_2 gnd vdd FILL
XFILL_85_DFFSR_184 gnd vdd FILL
XFILL_5_DFFSR_210 gnd vdd FILL
XFILL_85_DFFSR_195 gnd vdd FILL
XFILL_1_NOR2X1_190 gnd vdd FILL
XFILL_36_DFFSR_208 gnd vdd FILL
XFILL_5_DFFSR_221 gnd vdd FILL
XFILL_36_DFFSR_219 gnd vdd FILL
XFILL_5_DFFSR_232 gnd vdd FILL
XFILL_58_3 gnd vdd FILL
XFILL_5_DFFSR_243 gnd vdd FILL
XFILL_43_DFFSR_12 gnd vdd FILL
XFILL_5_DFFSR_254 gnd vdd FILL
XFILL_43_DFFSR_23 gnd vdd FILL
XFILL_5_DFFSR_265 gnd vdd FILL
XFILL_8_BUFX4_80 gnd vdd FILL
XFILL_8_BUFX4_91 gnd vdd FILL
XFILL_43_DFFSR_34 gnd vdd FILL
XFILL_14_NOR3X1_9 gnd vdd FILL
XFILL_43_DFFSR_45 gnd vdd FILL
XFILL_43_DFFSR_56 gnd vdd FILL
XFILL_63_DFFSR_108 gnd vdd FILL
XFILL_35_3_1 gnd vdd FILL
XFILL_43_DFFSR_67 gnd vdd FILL
XFILL_9_DFFSR_220 gnd vdd FILL
XFILL_43_DFFSR_78 gnd vdd FILL
XFILL_63_DFFSR_119 gnd vdd FILL
XFILL_9_DFFSR_231 gnd vdd FILL
XFILL_9_DFFSR_242 gnd vdd FILL
XFILL_43_DFFSR_89 gnd vdd FILL
XFILL_83_DFFSR_11 gnd vdd FILL
XFILL_10_NAND3X1_107 gnd vdd FILL
XFILL_9_DFFSR_253 gnd vdd FILL
XFILL_10_NAND3X1_118 gnd vdd FILL
XFILL_83_DFFSR_22 gnd vdd FILL
XFILL_9_DFFSR_264 gnd vdd FILL
XFILL_9_DFFSR_275 gnd vdd FILL
XFILL_10_NAND3X1_129 gnd vdd FILL
XFILL_83_DFFSR_33 gnd vdd FILL
XFILL_83_DFFSR_44 gnd vdd FILL
XFILL_67_DFFSR_107 gnd vdd FILL
XFILL_83_DFFSR_55 gnd vdd FILL
XFILL_12_DFFSR_11 gnd vdd FILL
XFILL_12_DFFSR_22 gnd vdd FILL
XFILL_83_DFFSR_66 gnd vdd FILL
XFILL_67_DFFSR_118 gnd vdd FILL
XFILL_1_MUX2X1_130 gnd vdd FILL
XFILL_83_DFFSR_77 gnd vdd FILL
XFILL_1_MUX2X1_141 gnd vdd FILL
XFILL_12_DFFSR_33 gnd vdd FILL
XFILL_83_DFFSR_88 gnd vdd FILL
XFILL_67_DFFSR_129 gnd vdd FILL
XFILL_1_MUX2X1_152 gnd vdd FILL
XFILL_12_DFFSR_44 gnd vdd FILL
XFILL_1_MUX2X1_163 gnd vdd FILL
XFILL_12_DFFSR_55 gnd vdd FILL
XFILL_83_DFFSR_99 gnd vdd FILL
XFILL_14_NAND3X1_16 gnd vdd FILL
XFILL_10_OAI21X1_8 gnd vdd FILL
XFILL_12_DFFSR_66 gnd vdd FILL
XFILL_14_NAND3X1_27 gnd vdd FILL
XFILL_1_MUX2X1_174 gnd vdd FILL
XFILL_12_DFFSR_77 gnd vdd FILL
XFILL_1_MUX2X1_185 gnd vdd FILL
XFILL_14_NAND3X1_38 gnd vdd FILL
XFILL_12_DFFSR_88 gnd vdd FILL
XFILL_14_NAND3X1_49 gnd vdd FILL
XFILL_12_DFFSR_99 gnd vdd FILL
XFILL_52_DFFSR_10 gnd vdd FILL
XFILL_52_DFFSR_21 gnd vdd FILL
XFILL_34_CLKBUF1_16 gnd vdd FILL
XFILL_52_DFFSR_32 gnd vdd FILL
XFILL_11_NOR2X1_10 gnd vdd FILL
XFILL_34_CLKBUF1_27 gnd vdd FILL
XFILL_52_DFFSR_43 gnd vdd FILL
XFILL_11_NOR2X1_21 gnd vdd FILL
XFILL_23_NOR3X1_7 gnd vdd FILL
XFILL_34_CLKBUF1_38 gnd vdd FILL
XFILL_21_DFFSR_230 gnd vdd FILL
XFILL_2_AOI22X1_4 gnd vdd FILL
XFILL_14_OAI21X1_7 gnd vdd FILL
XFILL_52_DFFSR_54 gnd vdd FILL
XFILL_11_NOR2X1_32 gnd vdd FILL
XFILL_11_NOR2X1_43 gnd vdd FILL
XFILL_21_DFFSR_241 gnd vdd FILL
XFILL_52_DFFSR_65 gnd vdd FILL
XFILL_52_DFFSR_76 gnd vdd FILL
XFILL_11_NOR2X1_54 gnd vdd FILL
XFILL_21_DFFSR_252 gnd vdd FILL
XFILL_11_NOR2X1_65 gnd vdd FILL
XFILL_52_DFFSR_87 gnd vdd FILL
XFILL_21_DFFSR_263 gnd vdd FILL
XFILL_21_DFFSR_274 gnd vdd FILL
XFILL_52_DFFSR_98 gnd vdd FILL
XFILL_11_NOR2X1_76 gnd vdd FILL
XFILL_2_INVX1_203 gnd vdd FILL
XFILL_9_MUX2X1_2 gnd vdd FILL
XFILL_2_INVX1_214 gnd vdd FILL
XFILL_11_NOR2X1_87 gnd vdd FILL
XFILL_1_DFFSR_5 gnd vdd FILL
XFILL_11_NOR2X1_98 gnd vdd FILL
XFILL_2_INVX1_225 gnd vdd FILL
XFILL_14_DFFSR_3 gnd vdd FILL
XFILL_6_AOI22X1_3 gnd vdd FILL
XFILL_25_DFFSR_240 gnd vdd FILL
XFILL_71_DFFSR_4 gnd vdd FILL
XFILL_21_DFFSR_20 gnd vdd FILL
XFILL_25_DFFSR_251 gnd vdd FILL
XFILL_21_DFFSR_31 gnd vdd FILL
XFILL_25_DFFSR_262 gnd vdd FILL
XFILL_21_DFFSR_42 gnd vdd FILL
XFILL_21_DFFSR_53 gnd vdd FILL
XFILL_25_DFFSR_273 gnd vdd FILL
XFILL_22_MUX2X1_18 gnd vdd FILL
XFILL_6_INVX1_202 gnd vdd FILL
XFILL_6_INVX1_213 gnd vdd FILL
XFILL_21_DFFSR_64 gnd vdd FILL
XFILL_22_MUX2X1_29 gnd vdd FILL
XFILL_21_DFFSR_75 gnd vdd FILL
XFILL_6_INVX1_224 gnd vdd FILL
XFILL_21_DFFSR_86 gnd vdd FILL
XFILL_21_DFFSR_97 gnd vdd FILL
XFILL_6_NOR3X1_8 gnd vdd FILL
XFILL_52_DFFSR_140 gnd vdd FILL
XFILL_52_DFFSR_151 gnd vdd FILL
XFILL_29_DFFSR_250 gnd vdd FILL
XFILL_52_DFFSR_162 gnd vdd FILL
XFILL_61_DFFSR_30 gnd vdd FILL
XFILL_52_DFFSR_173 gnd vdd FILL
XFILL_61_DFFSR_41 gnd vdd FILL
XFILL_29_DFFSR_261 gnd vdd FILL
XFILL_29_DFFSR_272 gnd vdd FILL
XFILL_61_DFFSR_52 gnd vdd FILL
XFILL_61_DFFSR_63 gnd vdd FILL
XFILL_52_DFFSR_184 gnd vdd FILL
XFILL_52_DFFSR_195 gnd vdd FILL
XFILL_4_NAND3X1_11 gnd vdd FILL
XFILL_61_DFFSR_74 gnd vdd FILL
XFILL_61_DFFSR_85 gnd vdd FILL
XFILL_4_NAND3X1_22 gnd vdd FILL
XFILL_61_DFFSR_96 gnd vdd FILL
XFILL_4_NAND3X1_33 gnd vdd FILL
XFILL_56_DFFSR_150 gnd vdd FILL
XFILL_4_NAND3X1_44 gnd vdd FILL
XFILL_26_3_1 gnd vdd FILL
XFILL_56_DFFSR_161 gnd vdd FILL
XFILL_4_NAND3X1_55 gnd vdd FILL
XFILL_1_3_1 gnd vdd FILL
XFILL_4_DFFSR_10 gnd vdd FILL
XFILL_4_DFFSR_21 gnd vdd FILL
XFILL_56_DFFSR_172 gnd vdd FILL
XFILL_8_NAND2X1_13 gnd vdd FILL
XFILL_4_NAND3X1_66 gnd vdd FILL
XFILL_8_NAND2X1_24 gnd vdd FILL
XFILL_4_DFFSR_32 gnd vdd FILL
XFILL_4_NAND3X1_77 gnd vdd FILL
XFILL_4_DFFSR_43 gnd vdd FILL
XFILL_56_DFFSR_183 gnd vdd FILL
XFILL_8_NAND2X1_35 gnd vdd FILL
XFILL_30_DFFSR_108 gnd vdd FILL
XFILL_4_NAND3X1_88 gnd vdd FILL
XFILL_56_DFFSR_194 gnd vdd FILL
XFILL_4_DFFSR_54 gnd vdd FILL
XFILL_36_DFFSR_7 gnd vdd FILL
XFILL_4_NAND3X1_99 gnd vdd FILL
XFILL_8_NAND2X1_46 gnd vdd FILL
XFILL_30_DFFSR_40 gnd vdd FILL
XFILL_8_NAND2X1_57 gnd vdd FILL
XFILL_4_DFFSR_65 gnd vdd FILL
XFILL_30_DFFSR_119 gnd vdd FILL
XFILL_4_DFFSR_76 gnd vdd FILL
XFILL_30_DFFSR_51 gnd vdd FILL
XFILL_8_NAND2X1_68 gnd vdd FILL
XFILL_8_NAND2X1_79 gnd vdd FILL
XFILL_4_DFFSR_87 gnd vdd FILL
XFILL_30_DFFSR_62 gnd vdd FILL
XFILL_4_DFFSR_98 gnd vdd FILL
XFILL_30_DFFSR_73 gnd vdd FILL
XFILL_30_DFFSR_84 gnd vdd FILL
XFILL_30_DFFSR_95 gnd vdd FILL
XFILL_34_DFFSR_107 gnd vdd FILL
XFILL_3_DFFSR_120 gnd vdd FILL
XFILL_34_DFFSR_118 gnd vdd FILL
XFILL_3_DFFSR_131 gnd vdd FILL
XFILL_11_NAND2X1_9 gnd vdd FILL
XFILL_3_DFFSR_142 gnd vdd FILL
XFILL_10_7_2 gnd vdd FILL
XFILL_34_DFFSR_129 gnd vdd FILL
XFILL_70_DFFSR_50 gnd vdd FILL
XFILL_3_DFFSR_153 gnd vdd FILL
XFILL_70_DFFSR_61 gnd vdd FILL
XFILL_11_AOI21X1_18 gnd vdd FILL
XFILL_70_DFFSR_72 gnd vdd FILL
XFILL_3_DFFSR_164 gnd vdd FILL
XFILL_70_DFFSR_83 gnd vdd FILL
XFILL_3_DFFSR_175 gnd vdd FILL
XFILL_11_AOI21X1_29 gnd vdd FILL
XFILL_3_DFFSR_186 gnd vdd FILL
XFILL_70_DFFSR_94 gnd vdd FILL
XFILL_3_DFFSR_197 gnd vdd FILL
XFILL_38_DFFSR_106 gnd vdd FILL
XFILL_7_DFFSR_130 gnd vdd FILL
XFILL_38_DFFSR_117 gnd vdd FILL
XFILL_38_DFFSR_128 gnd vdd FILL
XFILL_7_DFFSR_141 gnd vdd FILL
XFILL_7_DFFSR_152 gnd vdd FILL
XFILL_38_DFFSR_139 gnd vdd FILL
XFILL_11_MUX2X1_50 gnd vdd FILL
XFILL_7_DFFSR_163 gnd vdd FILL
XFILL_11_MUX2X1_61 gnd vdd FILL
XFILL_7_DFFSR_174 gnd vdd FILL
XFILL_10_NOR3X1_2 gnd vdd FILL
XFILL_11_MUX2X1_72 gnd vdd FILL
XFILL_11_MUX2X1_83 gnd vdd FILL
XFILL_8_AOI22X1_11 gnd vdd FILL
XFILL_7_DFFSR_185 gnd vdd FILL
XFILL_11_MUX2X1_94 gnd vdd FILL
XFILL_30_NOR3X1_19 gnd vdd FILL
XFILL_7_DFFSR_196 gnd vdd FILL
XFILL_9_4_1 gnd vdd FILL
XFILL_80_DFFSR_208 gnd vdd FILL
XFILL_80_DFFSR_219 gnd vdd FILL
XFILL_15_MUX2X1_60 gnd vdd FILL
XFILL_15_MUX2X1_71 gnd vdd FILL
XFILL_15_MUX2X1_82 gnd vdd FILL
XFILL_3_NOR3X1_20 gnd vdd FILL
XFILL_15_MUX2X1_93 gnd vdd FILL
XFILL_3_NOR3X1_31 gnd vdd FILL
XFILL_3_NOR3X1_42 gnd vdd FILL
XFILL_23_CLKBUF1_12 gnd vdd FILL
XFILL_23_CLKBUF1_23 gnd vdd FILL
XFILL_84_DFFSR_207 gnd vdd FILL
XFILL_23_CLKBUF1_34 gnd vdd FILL
XFILL_84_DFFSR_218 gnd vdd FILL
XFILL_84_DFFSR_229 gnd vdd FILL
XFILL_19_MUX2X1_70 gnd vdd FILL
XFILL_19_MUX2X1_81 gnd vdd FILL
XFILL_19_MUX2X1_92 gnd vdd FILL
XFILL_0_INVX1_102 gnd vdd FILL
XFILL_6_CLKBUF1_16 gnd vdd FILL
XFILL_7_NOR3X1_30 gnd vdd FILL
XFILL_0_INVX1_113 gnd vdd FILL
XFILL_6_CLKBUF1_27 gnd vdd FILL
XFILL_7_NOR3X1_41 gnd vdd FILL
XFILL_6_CLKBUF1_38 gnd vdd FILL
XFILL_7_NOR3X1_52 gnd vdd FILL
XFILL_0_INVX1_124 gnd vdd FILL
XFILL_17_3_1 gnd vdd FILL
XFILL_1_AOI21X1_13 gnd vdd FILL
XFILL_0_INVX1_135 gnd vdd FILL
XFILL_0_INVX1_146 gnd vdd FILL
XFILL_1_AOI21X1_24 gnd vdd FILL
XFILL_0_INVX1_157 gnd vdd FILL
XFILL_1_AOI21X1_35 gnd vdd FILL
XFILL_0_INVX1_168 gnd vdd FILL
XFILL_23_DFFSR_150 gnd vdd FILL
XFILL_23_DFFSR_161 gnd vdd FILL
XFILL_1_AOI21X1_46 gnd vdd FILL
XFILL_23_DFFSR_172 gnd vdd FILL
XFILL_11_OAI22X1_15 gnd vdd FILL
XFILL_0_INVX1_179 gnd vdd FILL
XFILL_1_AOI21X1_57 gnd vdd FILL
XFILL_60_6_2 gnd vdd FILL
XFILL_1_AOI21X1_68 gnd vdd FILL
XFILL_4_INVX1_101 gnd vdd FILL
XFILL_4_INVX1_112 gnd vdd FILL
XFILL_23_DFFSR_183 gnd vdd FILL
XFILL_11_OAI22X1_26 gnd vdd FILL
XFILL_1_AOI21X1_79 gnd vdd FILL
XFILL_4_INVX1_123 gnd vdd FILL
XFILL_23_DFFSR_194 gnd vdd FILL
XFILL_11_OAI22X1_37 gnd vdd FILL
XFILL_4_NOR2X1_101 gnd vdd FILL
XFILL_11_OAI22X1_48 gnd vdd FILL
XFILL_4_INVX1_134 gnd vdd FILL
XFILL_4_NOR2X1_112 gnd vdd FILL
XFILL_15_OAI21X1_17 gnd vdd FILL
XFILL_4_NOR2X1_123 gnd vdd FILL
XFILL_4_INVX1_145 gnd vdd FILL
XFILL_4_INVX1_156 gnd vdd FILL
XFILL_15_OAI21X1_28 gnd vdd FILL
XFILL_4_INVX1_167 gnd vdd FILL
XFILL_4_NOR2X1_134 gnd vdd FILL
XFILL_15_OAI21X1_39 gnd vdd FILL
XFILL_27_DFFSR_160 gnd vdd FILL
XFILL_4_NOR2X1_145 gnd vdd FILL
XFILL_4_NOR2X1_156 gnd vdd FILL
XFILL_27_DFFSR_171 gnd vdd FILL
XFILL_4_INVX1_178 gnd vdd FILL
XFILL_4_INVX1_189 gnd vdd FILL
XFILL_4_NOR2X1_167 gnd vdd FILL
XFILL_27_DFFSR_182 gnd vdd FILL
XFILL_4_NOR2X1_178 gnd vdd FILL
XFILL_27_DFFSR_193 gnd vdd FILL
XFILL_11_INVX8_1 gnd vdd FILL
XFILL_4_NOR2X1_189 gnd vdd FILL
XFILL_10_NAND3X1_80 gnd vdd FILL
XFILL_2_NOR3X1_1 gnd vdd FILL
XFILL_10_NAND3X1_91 gnd vdd FILL
XFILL_23_NOR3X1_50 gnd vdd FILL
XFILL_21_MUX2X1_103 gnd vdd FILL
XFILL_21_MUX2X1_114 gnd vdd FILL
XFILL_21_MUX2X1_125 gnd vdd FILL
XFILL_2_OAI22X1_7 gnd vdd FILL
XFILL_21_MUX2X1_136 gnd vdd FILL
XFILL_21_MUX2X1_147 gnd vdd FILL
XFILL_21_MUX2X1_158 gnd vdd FILL
XFILL_73_DFFSR_250 gnd vdd FILL
XFILL_21_MUX2X1_169 gnd vdd FILL
XFILL_53_DFFSR_1 gnd vdd FILL
XFILL_73_DFFSR_261 gnd vdd FILL
XFILL_73_DFFSR_272 gnd vdd FILL
XFILL_4_MUX2X1_107 gnd vdd FILL
XFILL_4_MUX2X1_118 gnd vdd FILL
XFILL_0_DFFSR_80 gnd vdd FILL
XFILL_4_MUX2X1_129 gnd vdd FILL
XFILL_0_DFFSR_91 gnd vdd FILL
XFILL_9_NOR2X1_201 gnd vdd FILL
XFILL_6_OAI22X1_6 gnd vdd FILL
XFILL_1_OAI22X1_10 gnd vdd FILL
XFILL_1_OAI22X1_21 gnd vdd FILL
XFILL_63_1 gnd vdd FILL
XFILL_1_OAI22X1_32 gnd vdd FILL
XFILL_1_OAI22X1_43 gnd vdd FILL
XFILL_77_DFFSR_260 gnd vdd FILL
XFILL_77_DFFSR_271 gnd vdd FILL
XFILL_32_CLKBUF1_1 gnd vdd FILL
XFILL_5_OAI21X1_12 gnd vdd FILL
XFILL_5_OAI21X1_23 gnd vdd FILL
XFILL_51_DFFSR_207 gnd vdd FILL
XFILL_5_OAI21X1_34 gnd vdd FILL
XFILL_51_DFFSR_218 gnd vdd FILL
XFILL_5_OAI21X1_45 gnd vdd FILL
XFILL_51_DFFSR_229 gnd vdd FILL
XFILL_5_DFFSR_6 gnd vdd FILL
XFILL_55_DFFSR_206 gnd vdd FILL
XFILL_18_DFFSR_4 gnd vdd FILL
XFILL_55_DFFSR_217 gnd vdd FILL
XFILL_51_6_2 gnd vdd FILL
XFILL_55_DFFSR_228 gnd vdd FILL
XFILL_75_DFFSR_5 gnd vdd FILL
XFILL_55_DFFSR_239 gnd vdd FILL
XFILL_50_1_1 gnd vdd FILL
XFILL_11_NAND3X1_108 gnd vdd FILL
XFILL_9_BUFX4_14 gnd vdd FILL
XFILL_9_BUFX4_25 gnd vdd FILL
XFILL_11_NAND3X1_119 gnd vdd FILL
XFILL_9_BUFX4_36 gnd vdd FILL
XFILL_9_BUFX4_47 gnd vdd FILL
XFILL_82_DFFSR_106 gnd vdd FILL
XFILL_9_BUFX4_58 gnd vdd FILL
XFILL_12_CLKBUF1_30 gnd vdd FILL
XFILL_59_DFFSR_205 gnd vdd FILL
XFILL_9_BUFX4_69 gnd vdd FILL
XFILL_82_DFFSR_117 gnd vdd FILL
XFILL_59_DFFSR_216 gnd vdd FILL
XFILL_12_CLKBUF1_41 gnd vdd FILL
XFILL_59_DFFSR_227 gnd vdd FILL
XFILL_82_DFFSR_128 gnd vdd FILL
XFILL_59_DFFSR_238 gnd vdd FILL
XFILL_82_DFFSR_139 gnd vdd FILL
XFILL_59_DFFSR_249 gnd vdd FILL
XFILL_86_DFFSR_105 gnd vdd FILL
XFILL_2_DFFSR_209 gnd vdd FILL
XFILL_86_DFFSR_116 gnd vdd FILL
XFILL_86_DFFSR_127 gnd vdd FILL
XFILL_86_DFFSR_138 gnd vdd FILL
XFILL_86_DFFSR_149 gnd vdd FILL
XFILL_6_DFFSR_208 gnd vdd FILL
XFILL_3_NAND3X1_8 gnd vdd FILL
XFILL_6_DFFSR_219 gnd vdd FILL
XFILL_10_NOR2X1_170 gnd vdd FILL
XFILL_10_NOR2X1_181 gnd vdd FILL
XFILL_10_NOR2X1_192 gnd vdd FILL
XFILL_40_DFFSR_250 gnd vdd FILL
XFILL_59_7_2 gnd vdd FILL
XFILL_40_DFFSR_261 gnd vdd FILL
XFILL_40_DFFSR_272 gnd vdd FILL
XFILL_7_NAND3X1_7 gnd vdd FILL
XFILL_58_2_1 gnd vdd FILL
XFILL_44_DFFSR_260 gnd vdd FILL
XFILL_44_DFFSR_271 gnd vdd FILL
XFILL_13_BUFX4_30 gnd vdd FILL
XFILL_12_BUFX4_4 gnd vdd FILL
XFILL_13_BUFX4_41 gnd vdd FILL
XFILL_10_MUX2X1_110 gnd vdd FILL
XFILL_13_BUFX4_52 gnd vdd FILL
XFILL_10_MUX2X1_121 gnd vdd FILL
XFILL_13_BUFX4_63 gnd vdd FILL
XFILL_13_BUFX4_74 gnd vdd FILL
XFILL_10_MUX2X1_132 gnd vdd FILL
XFILL_13_BUFX4_85 gnd vdd FILL
XFILL_10_MUX2X1_143 gnd vdd FILL
XFILL_71_DFFSR_160 gnd vdd FILL
XFILL_13_BUFX4_96 gnd vdd FILL
XFILL_10_MUX2X1_154 gnd vdd FILL
XFILL_10_MUX2X1_165 gnd vdd FILL
XFILL_71_DFFSR_171 gnd vdd FILL
XFILL_48_DFFSR_270 gnd vdd FILL
XFILL_42_6_2 gnd vdd FILL
XFILL_10_MUX2X1_176 gnd vdd FILL
XFILL_71_DFFSR_182 gnd vdd FILL
XFILL_62_DFFSR_19 gnd vdd FILL
XFILL_10_MUX2X1_187 gnd vdd FILL
XFILL_71_DFFSR_193 gnd vdd FILL
XFILL_22_DFFSR_206 gnd vdd FILL
XFILL_41_1_1 gnd vdd FILL
XFILL_22_DFFSR_217 gnd vdd FILL
XFILL_22_DFFSR_228 gnd vdd FILL
XFILL_22_DFFSR_239 gnd vdd FILL
XFILL_75_DFFSR_170 gnd vdd FILL
XFILL_75_DFFSR_181 gnd vdd FILL
XFILL_75_DFFSR_192 gnd vdd FILL
XFILL_26_DFFSR_205 gnd vdd FILL
XAOI22X1_4 NOR2X1_40/Y INVX1_175/A INVX1_170/A NOR2X1_41/Y gnd AOI22X1_4/Y vdd AOI22X1
XFILL_26_DFFSR_216 gnd vdd FILL
XFILL_26_DFFSR_227 gnd vdd FILL
XFILL_26_DFFSR_238 gnd vdd FILL
XFILL_31_DFFSR_18 gnd vdd FILL
XFILL_26_DFFSR_249 gnd vdd FILL
XFILL_31_DFFSR_29 gnd vdd FILL
XFILL_7_INVX1_20 gnd vdd FILL
XFILL_7_INVX1_31 gnd vdd FILL
XINVX1_203 DFFSR_87/Q gnd INVX1_203/Y vdd INVX1
XFILL_79_DFFSR_180 gnd vdd FILL
XFILL_7_INVX1_42 gnd vdd FILL
XFILL_7_INVX1_53 gnd vdd FILL
XINVX1_214 DFFSR_75/Q gnd INVX1_214/Y vdd INVX1
XFILL_79_DFFSR_191 gnd vdd FILL
XFILL_8_AND2X2_1 gnd vdd FILL
XFILL_53_DFFSR_105 gnd vdd FILL
XINVX1_225 DFFSR_60/Q gnd OAI22X1_9/C vdd INVX1
XFILL_7_INVX1_64 gnd vdd FILL
XFILL_53_DFFSR_116 gnd vdd FILL
XFILL_7_INVX1_75 gnd vdd FILL
XFILL_7_INVX1_86 gnd vdd FILL
XFILL_53_DFFSR_127 gnd vdd FILL
XFILL_53_DFFSR_138 gnd vdd FILL
XFILL_7_INVX1_97 gnd vdd FILL
XFILL_71_DFFSR_17 gnd vdd FILL
XFILL_53_DFFSR_149 gnd vdd FILL
XFILL_71_DFFSR_28 gnd vdd FILL
XFILL_71_DFFSR_39 gnd vdd FILL
XFILL_14_MUX2X1_7 gnd vdd FILL
XFILL_57_DFFSR_104 gnd vdd FILL
XFILL_57_DFFSR_115 gnd vdd FILL
XFILL_57_DFFSR_126 gnd vdd FILL
XFILL_57_DFFSR_137 gnd vdd FILL
XFILL_57_DFFSR_148 gnd vdd FILL
XNAND2X1_14 INVX2_1/A INVX1_3/A gnd MUX2X1_95/S vdd NAND2X1
XFILL_0_MUX2X1_160 gnd vdd FILL
XFILL_13_NAND3X1_13 gnd vdd FILL
XFILL_5_BUFX4_40 gnd vdd FILL
XFILL_0_MUX2X1_171 gnd vdd FILL
XFILL_57_DFFSR_159 gnd vdd FILL
XNAND2X1_25 AND2X2_5/B AND2X2_6/A gnd NOR2X1_40/B vdd NAND2X1
XFILL_13_NAND3X1_24 gnd vdd FILL
XFILL_49_2_1 gnd vdd FILL
XFILL_0_MUX2X1_182 gnd vdd FILL
XNAND2X1_36 BUFX4_103/Y NOR2X1_31/Y gnd OAI22X1_50/B vdd NAND2X1
XFILL_13_NAND3X1_35 gnd vdd FILL
XFILL_2_INVX8_4 gnd vdd FILL
XFILL_5_BUFX4_51 gnd vdd FILL
XFILL_13_NAND3X1_46 gnd vdd FILL
XFILL_0_MUX2X1_193 gnd vdd FILL
XFILL_0_DFFSR_108 gnd vdd FILL
XFILL_40_DFFSR_16 gnd vdd FILL
XFILL_5_BUFX4_62 gnd vdd FILL
XNAND2X1_47 AND2X2_3/B AND2X2_6/A gnd NOR3X1_5/C vdd NAND2X1
XFILL_13_NAND3X1_57 gnd vdd FILL
XFILL_5_BUFX4_73 gnd vdd FILL
XNAND2X1_58 BUFX4_102/Y NOR2X1_38/Y gnd OAI21X1_6/B vdd NAND2X1
XFILL_40_DFFSR_27 gnd vdd FILL
XFILL_5_BUFX4_84 gnd vdd FILL
XFILL_15_INVX8_2 gnd vdd FILL
XFILL_13_NAND3X1_68 gnd vdd FILL
XNAND2X1_69 NAND2X1_69/A NAND2X1_69/B gnd NOR3X1_31/A vdd NAND2X1
XFILL_0_DFFSR_119 gnd vdd FILL
XFILL_33_CLKBUF1_13 gnd vdd FILL
XFILL_5_BUFX4_95 gnd vdd FILL
XFILL_33_CLKBUF1_24 gnd vdd FILL
XFILL_40_DFFSR_38 gnd vdd FILL
XFILL_13_NAND3X1_79 gnd vdd FILL
XFILL_33_CLKBUF1_35 gnd vdd FILL
XFILL_40_DFFSR_49 gnd vdd FILL
XFILL_11_DFFSR_260 gnd vdd FILL
XFILL_4_DFFSR_107 gnd vdd FILL
XFILL_11_DFFSR_271 gnd vdd FILL
XFILL_80_DFFSR_15 gnd vdd FILL
XFILL_80_DFFSR_26 gnd vdd FILL
XFILL_4_DFFSR_118 gnd vdd FILL
XFILL_80_DFFSR_37 gnd vdd FILL
XFILL_4_DFFSR_129 gnd vdd FILL
XFILL_23_MUX2X1_5 gnd vdd FILL
XFILL_80_DFFSR_48 gnd vdd FILL
XFILL_80_DFFSR_59 gnd vdd FILL
XFILL_33_6_2 gnd vdd FILL
XFILL_28_4 gnd vdd FILL
XFILL_32_1_1 gnd vdd FILL
XFILL_8_DFFSR_106 gnd vdd FILL
XFILL_15_DFFSR_270 gnd vdd FILL
XFILL_57_DFFSR_2 gnd vdd FILL
XFILL_8_DFFSR_117 gnd vdd FILL
XFILL_12_MUX2X1_15 gnd vdd FILL
XFILL_7_NOR2X1_8 gnd vdd FILL
XFILL_8_DFFSR_128 gnd vdd FILL
XFILL_12_MUX2X1_26 gnd vdd FILL
XFILL_12_MUX2X1_37 gnd vdd FILL
XFILL_8_DFFSR_139 gnd vdd FILL
XFILL_3_AOI21X1_2 gnd vdd FILL
XFILL_12_MUX2X1_48 gnd vdd FILL
XFILL_12_MUX2X1_59 gnd vdd FILL
XFILL_42_DFFSR_170 gnd vdd FILL
XFILL_0_NOR3X1_19 gnd vdd FILL
XFILL_16_MUX2X1_14 gnd vdd FILL
XFILL_42_DFFSR_181 gnd vdd FILL
XFILL_16_MUX2X1_25 gnd vdd FILL
XFILL_42_DFFSR_192 gnd vdd FILL
XFILL_16_MUX2X1_36 gnd vdd FILL
XFILL_16_MUX2X1_47 gnd vdd FILL
XFILL_7_AOI21X1_1 gnd vdd FILL
XFILL_16_MUX2X1_58 gnd vdd FILL
XFILL_3_NAND3X1_30 gnd vdd FILL
XFILL_6_MUX2X1_6 gnd vdd FILL
XFILL_16_MUX2X1_69 gnd vdd FILL
XNOR3X1_2 NOR3X1_9/A NOR3X1_9/B NOR3X1_2/C gnd NOR3X1_2/Y vdd NOR3X1
XFILL_3_NAND3X1_41 gnd vdd FILL
XFILL_3_NAND3X1_52 gnd vdd FILL
XFILL_7_NAND2X1_10 gnd vdd FILL
XFILL_4_NOR3X1_18 gnd vdd FILL
XFILL_3_NAND3X1_63 gnd vdd FILL
XFILL_46_DFFSR_180 gnd vdd FILL
XFILL_4_NOR3X1_29 gnd vdd FILL
XFILL_7_NAND2X1_21 gnd vdd FILL
XFILL_3_NAND3X1_74 gnd vdd FILL
XFILL_41_DFFSR_8 gnd vdd FILL
XFILL_7_NAND2X1_32 gnd vdd FILL
XFILL_20_DFFSR_105 gnd vdd FILL
XFILL_3_NAND3X1_85 gnd vdd FILL
XFILL_46_DFFSR_191 gnd vdd FILL
XFILL_7_NAND2X1_43 gnd vdd FILL
XFILL_9_DFFSR_7 gnd vdd FILL
XFILL_3_NAND3X1_96 gnd vdd FILL
XFILL_20_DFFSR_116 gnd vdd FILL
XFILL_7_NAND2X1_54 gnd vdd FILL
XFILL_7_NAND2X1_65 gnd vdd FILL
XFILL_20_DFFSR_127 gnd vdd FILL
XFILL_20_DFFSR_138 gnd vdd FILL
XFILL_7_NAND2X1_76 gnd vdd FILL
XFILL_20_DFFSR_149 gnd vdd FILL
XFILL_79_DFFSR_6 gnd vdd FILL
XFILL_7_NAND2X1_87 gnd vdd FILL
XFILL_8_NOR3X1_17 gnd vdd FILL
XFILL_8_NOR3X1_28 gnd vdd FILL
XFILL_8_NOR3X1_39 gnd vdd FILL
XFILL_24_DFFSR_104 gnd vdd FILL
XFILL_15_CLKBUF1_18 gnd vdd FILL
XFILL_24_DFFSR_115 gnd vdd FILL
XFILL_15_CLKBUF1_29 gnd vdd FILL
XFILL_24_DFFSR_126 gnd vdd FILL
XFILL_24_DFFSR_137 gnd vdd FILL
XFILL_24_DFFSR_148 gnd vdd FILL
XFILL_10_AOI21X1_15 gnd vdd FILL
XFILL_10_AOI21X1_26 gnd vdd FILL
XFILL_24_DFFSR_159 gnd vdd FILL
XFILL_10_AOI21X1_37 gnd vdd FILL
XFILL_10_AOI21X1_48 gnd vdd FILL
XFILL_10_AOI21X1_59 gnd vdd FILL
XFILL_28_DFFSR_103 gnd vdd FILL
XFILL_1_DFFSR_14 gnd vdd FILL
XFILL_11_NOR2X1_2 gnd vdd FILL
XFILL_28_DFFSR_114 gnd vdd FILL
XFILL_1_DFFSR_25 gnd vdd FILL
XFILL_1_DFFSR_36 gnd vdd FILL
XFILL_28_DFFSR_125 gnd vdd FILL
XFILL_1_DFFSR_47 gnd vdd FILL
XFILL_28_DFFSR_136 gnd vdd FILL
XFILL_1_DFFSR_58 gnd vdd FILL
XFILL_28_DFFSR_147 gnd vdd FILL
XFILL_28_DFFSR_158 gnd vdd FILL
XFILL_1_DFFSR_69 gnd vdd FILL
XFILL_28_DFFSR_169 gnd vdd FILL
XFILL_20_NOR3X1_16 gnd vdd FILL
XFILL_24_6_2 gnd vdd FILL
XFILL_20_NOR3X1_27 gnd vdd FILL
XFILL_20_NOR3X1_38 gnd vdd FILL
XFILL_20_NOR3X1_49 gnd vdd FILL
XFILL_3_INVX1_90 gnd vdd FILL
XFILL_23_1_1 gnd vdd FILL
XFILL_70_DFFSR_205 gnd vdd FILL
XFILL_3_BUFX2_10 gnd vdd FILL
XFILL_70_DFFSR_216 gnd vdd FILL
XFILL_70_DFFSR_227 gnd vdd FILL
XFILL_70_DFFSR_238 gnd vdd FILL
XFILL_49_DFFSR_60 gnd vdd FILL
XFILL_49_DFFSR_71 gnd vdd FILL
XFILL_12_NAND3X1_109 gnd vdd FILL
XFILL_49_DFFSR_82 gnd vdd FILL
XFILL_70_DFFSR_249 gnd vdd FILL
XFILL_49_DFFSR_93 gnd vdd FILL
XFILL_24_NOR3X1_15 gnd vdd FILL
XFILL_24_NOR3X1_26 gnd vdd FILL
XFILL_24_NOR3X1_37 gnd vdd FILL
XFILL_22_CLKBUF1_20 gnd vdd FILL
XFILL_24_NOR3X1_48 gnd vdd FILL
XFILL_22_CLKBUF1_31 gnd vdd FILL
XFILL_74_DFFSR_204 gnd vdd FILL
XFILL_74_DFFSR_215 gnd vdd FILL
XFILL_22_CLKBUF1_42 gnd vdd FILL
XFILL_74_DFFSR_226 gnd vdd FILL
XFILL_74_DFFSR_237 gnd vdd FILL
XFILL_74_DFFSR_248 gnd vdd FILL
XFILL_28_NOR3X1_14 gnd vdd FILL
XFILL_5_CLKBUF1_13 gnd vdd FILL
XFILL_74_DFFSR_259 gnd vdd FILL
XFILL_3_BUFX4_7 gnd vdd FILL
XFILL_5_CLKBUF1_24 gnd vdd FILL
XFILL_28_NOR3X1_25 gnd vdd FILL
XFILL_28_NOR3X1_36 gnd vdd FILL
XFILL_5_CLKBUF1_35 gnd vdd FILL
XFILL_28_NOR3X1_47 gnd vdd FILL
XFILL_78_DFFSR_203 gnd vdd FILL
XFILL_18_DFFSR_70 gnd vdd FILL
XFILL_13_MUX2X1_109 gnd vdd FILL
XOAI22X1_7 OAI22X1_7/A OAI22X1_7/B OAI22X1_7/C OAI22X1_7/D gnd OAI22X1_7/Y vdd OAI22X1
XFILL_0_AOI21X1_10 gnd vdd FILL
XFILL_18_DFFSR_81 gnd vdd FILL
XFILL_18_DFFSR_92 gnd vdd FILL
XFILL_0_AOI21X1_21 gnd vdd FILL
XFILL_78_DFFSR_214 gnd vdd FILL
XFILL_0_AOI21X1_32 gnd vdd FILL
XFILL_78_DFFSR_225 gnd vdd FILL
XFILL_0_AOI21X1_43 gnd vdd FILL
XFILL_78_DFFSR_236 gnd vdd FILL
XFILL_78_DFFSR_247 gnd vdd FILL
XFILL_2_CLKBUF1_1 gnd vdd FILL
XFILL_0_AOI21X1_54 gnd vdd FILL
XFILL_10_OAI22X1_12 gnd vdd FILL
XFILL_13_DFFSR_180 gnd vdd FILL
XFILL_10_OAI22X1_23 gnd vdd FILL
XFILL_78_DFFSR_258 gnd vdd FILL
XFILL_0_AOI21X1_65 gnd vdd FILL
XFILL_78_DFFSR_269 gnd vdd FILL
XFILL_0_AOI21X1_76 gnd vdd FILL
XFILL_10_OAI22X1_34 gnd vdd FILL
XFILL_13_DFFSR_191 gnd vdd FILL
XFILL_10_OAI22X1_45 gnd vdd FILL
XFILL_58_DFFSR_80 gnd vdd FILL
XFILL_14_OAI21X1_14 gnd vdd FILL
XFILL_58_DFFSR_91 gnd vdd FILL
XFILL_3_NOR2X1_120 gnd vdd FILL
XFILL_14_OAI21X1_25 gnd vdd FILL
XFILL_3_NOR2X1_131 gnd vdd FILL
XFILL_7_7_2 gnd vdd FILL
XFILL_14_OAI21X1_36 gnd vdd FILL
XFILL_14_OAI21X1_47 gnd vdd FILL
XFILL_3_NOR2X1_142 gnd vdd FILL
XFILL_3_NOR2X1_153 gnd vdd FILL
XFILL_3_NOR2X1_1 gnd vdd FILL
XFILL_6_2_1 gnd vdd FILL
XFILL_3_NOR2X1_164 gnd vdd FILL
XFILL_17_DFFSR_190 gnd vdd FILL
XFILL_3_NOR2X1_175 gnd vdd FILL
XFILL_3_NOR2X1_186 gnd vdd FILL
XFILL_3_NOR2X1_197 gnd vdd FILL
XFILL_27_DFFSR_90 gnd vdd FILL
XFILL_20_MUX2X1_100 gnd vdd FILL
XFILL_20_MUX2X1_111 gnd vdd FILL
XFILL_20_MUX2X1_122 gnd vdd FILL
XFILL_15_6_2 gnd vdd FILL
XFILL_20_MUX2X1_133 gnd vdd FILL
XFILL_20_MUX2X1_144 gnd vdd FILL
XFILL_20_MUX2X1_155 gnd vdd FILL
XFILL_14_1_1 gnd vdd FILL
XFILL_20_MUX2X1_166 gnd vdd FILL
XFILL_3_MUX2X1_104 gnd vdd FILL
XFILL_20_MUX2X1_177 gnd vdd FILL
XFILL_3_MUX2X1_115 gnd vdd FILL
XFILL_20_MUX2X1_188 gnd vdd FILL
XFILL_3_MUX2X1_126 gnd vdd FILL
XFILL_3_MUX2X1_137 gnd vdd FILL
XFILL_3_MUX2X1_148 gnd vdd FILL
XFILL_14_BUFX4_19 gnd vdd FILL
XFILL_3_MUX2X1_159 gnd vdd FILL
XFILL_0_OAI22X1_40 gnd vdd FILL
XFILL_0_OAI22X1_51 gnd vdd FILL
XDFFSR_209 INVX1_85/A DFFSR_57/CLK DFFSR_90/R vdd MUX2X1_72/Y gnd vdd DFFSR
XFILL_4_OAI21X1_20 gnd vdd FILL
XFILL_19_INVX8_3 gnd vdd FILL
XFILL_4_OAI21X1_31 gnd vdd FILL
XFILL_41_DFFSR_204 gnd vdd FILL
XFILL_41_DFFSR_215 gnd vdd FILL
XFILL_0_NOR2X1_30 gnd vdd FILL
XFILL_4_OAI21X1_42 gnd vdd FILL
XFILL_3_OAI21X1_5 gnd vdd FILL
XFILL_41_DFFSR_226 gnd vdd FILL
XFILL_0_NOR2X1_41 gnd vdd FILL
XFILL_41_DFFSR_237 gnd vdd FILL
XFILL_0_NOR2X1_52 gnd vdd FILL
XFILL_41_DFFSR_248 gnd vdd FILL
XFILL_0_NOR2X1_63 gnd vdd FILL
XFILL_0_NOR2X1_74 gnd vdd FILL
XFILL_41_DFFSR_259 gnd vdd FILL
XFILL_0_NOR2X1_85 gnd vdd FILL
XFILL_0_NOR2X1_96 gnd vdd FILL
XFILL_23_DFFSR_5 gnd vdd FILL
XFILL_45_DFFSR_203 gnd vdd FILL
XFILL_45_DFFSR_214 gnd vdd FILL
XFILL_7_OAI21X1_4 gnd vdd FILL
XFILL_45_DFFSR_225 gnd vdd FILL
XFILL_4_NOR2X1_40 gnd vdd FILL
XFILL_80_DFFSR_6 gnd vdd FILL
XFILL_45_DFFSR_236 gnd vdd FILL
XFILL_4_NOR2X1_51 gnd vdd FILL
XFILL_45_DFFSR_247 gnd vdd FILL
XFILL_4_NOR2X1_62 gnd vdd FILL
XFILL_45_DFFSR_258 gnd vdd FILL
XFILL_4_NOR2X1_73 gnd vdd FILL
XFILL_45_DFFSR_269 gnd vdd FILL
XFILL_4_NOR2X1_84 gnd vdd FILL
XFILL_49_DFFSR_202 gnd vdd FILL
XFILL_4_NOR2X1_95 gnd vdd FILL
XFILL_72_DFFSR_103 gnd vdd FILL
XFILL_72_DFFSR_114 gnd vdd FILL
XFILL_49_DFFSR_213 gnd vdd FILL
XFILL_72_DFFSR_125 gnd vdd FILL
XFILL_49_DFFSR_224 gnd vdd FILL
XFILL_72_DFFSR_136 gnd vdd FILL
XFILL_49_DFFSR_235 gnd vdd FILL
XFILL_8_NOR2X1_50 gnd vdd FILL
XFILL_12_OAI22X1_1 gnd vdd FILL
XFILL_49_DFFSR_246 gnd vdd FILL
XFILL_72_DFFSR_147 gnd vdd FILL
XFILL_72_DFFSR_158 gnd vdd FILL
XFILL_8_NOR2X1_61 gnd vdd FILL
XFILL_49_DFFSR_257 gnd vdd FILL
XFILL_72_DFFSR_169 gnd vdd FILL
XFILL_8_NOR2X1_72 gnd vdd FILL
XFILL_49_DFFSR_268 gnd vdd FILL
XFILL_8_NOR2X1_83 gnd vdd FILL
XFILL_65_5_2 gnd vdd FILL
XFILL_8_NOR2X1_94 gnd vdd FILL
XFILL_76_DFFSR_102 gnd vdd FILL
XFILL_76_DFFSR_113 gnd vdd FILL
XFILL_76_DFFSR_124 gnd vdd FILL
XFILL_64_0_1 gnd vdd FILL
XFILL_6_NAND3X1_18 gnd vdd FILL
XFILL_76_DFFSR_135 gnd vdd FILL
XFILL_6_NAND3X1_29 gnd vdd FILL
XFILL_76_DFFSR_146 gnd vdd FILL
XFILL_76_DFFSR_157 gnd vdd FILL
XFILL_76_DFFSR_168 gnd vdd FILL
XFILL_76_DFFSR_179 gnd vdd FILL
XFILL_45_DFFSR_9 gnd vdd FILL
XFILL_6_BUFX4_18 gnd vdd FILL
XFILL_6_BUFX4_29 gnd vdd FILL
XFILL_26_1 gnd vdd FILL
XFILL_0_NAND2X1_7 gnd vdd FILL
XFILL_4_NAND2X1_6 gnd vdd FILL
XFILL_0_MUX2X1_70 gnd vdd FILL
XFILL_0_MUX2X1_81 gnd vdd FILL
XFILL_13_AND2X2_6 gnd vdd FILL
XFILL_0_MUX2X1_92 gnd vdd FILL
XFILL_8_NAND2X1_5 gnd vdd FILL
XFILL_61_DFFSR_190 gnd vdd FILL
XFILL_12_DFFSR_203 gnd vdd FILL
XFILL_12_DFFSR_214 gnd vdd FILL
XFILL_12_DFFSR_225 gnd vdd FILL
XFILL_12_DFFSR_236 gnd vdd FILL
XFILL_4_MUX2X1_80 gnd vdd FILL
XFILL_4_MUX2X1_91 gnd vdd FILL
XFILL_12_DFFSR_247 gnd vdd FILL
XFILL_12_DFFSR_258 gnd vdd FILL
XFILL_12_DFFSR_269 gnd vdd FILL
XFILL_10_BUFX4_12 gnd vdd FILL
XFILL_16_DFFSR_202 gnd vdd FILL
XFILL_25_CLKBUF1_19 gnd vdd FILL
XFILL_10_BUFX4_23 gnd vdd FILL
XFILL_13_NAND3X1_2 gnd vdd FILL
XFILL_16_DFFSR_213 gnd vdd FILL
XFILL_16_DFFSR_224 gnd vdd FILL
XFILL_10_BUFX4_34 gnd vdd FILL
XFILL_10_BUFX4_45 gnd vdd FILL
XFILL_56_5_2 gnd vdd FILL
XFILL_16_DFFSR_235 gnd vdd FILL
XFILL_10_BUFX4_56 gnd vdd FILL
XFILL_16_DFFSR_246 gnd vdd FILL
XFILL_8_MUX2X1_90 gnd vdd FILL
XFILL_10_BUFX4_67 gnd vdd FILL
XFILL_55_0_1 gnd vdd FILL
XFILL_10_BUFX4_78 gnd vdd FILL
XFILL_7_BUFX4_8 gnd vdd FILL
XFILL_16_DFFSR_257 gnd vdd FILL
XFILL_16_DFFSR_268 gnd vdd FILL
XFILL_10_BUFX4_89 gnd vdd FILL
XFILL_43_DFFSR_102 gnd vdd FILL
XFILL_43_DFFSR_113 gnd vdd FILL
XFILL_43_DFFSR_124 gnd vdd FILL
XFILL_43_DFFSR_135 gnd vdd FILL
XFILL_43_DFFSR_146 gnd vdd FILL
XFILL_43_DFFSR_157 gnd vdd FILL
XFILL_43_DFFSR_168 gnd vdd FILL
XFILL_43_DFFSR_179 gnd vdd FILL
XFILL_47_DFFSR_101 gnd vdd FILL
XFILL_47_DFFSR_112 gnd vdd FILL
XFILL_6_NOR2X1_108 gnd vdd FILL
XFILL_47_DFFSR_123 gnd vdd FILL
XFILL_47_DFFSR_134 gnd vdd FILL
XFILL_6_NOR2X1_119 gnd vdd FILL
XFILL_47_DFFSR_145 gnd vdd FILL
XFILL_12_NAND3X1_10 gnd vdd FILL
XFILL_47_DFFSR_156 gnd vdd FILL
XFILL_12_NAND3X1_21 gnd vdd FILL
XFILL_47_DFFSR_167 gnd vdd FILL
XFILL_12_NAND3X1_32 gnd vdd FILL
XFILL_47_DFFSR_178 gnd vdd FILL
XFILL_12_NAND3X1_43 gnd vdd FILL
XFILL_4_INVX1_13 gnd vdd FILL
XFILL_47_DFFSR_189 gnd vdd FILL
XFILL_12_NAND3X1_54 gnd vdd FILL
XFILL_4_INVX1_24 gnd vdd FILL
XFILL_12_NAND3X1_65 gnd vdd FILL
XFILL_4_INVX1_35 gnd vdd FILL
XFILL_32_CLKBUF1_10 gnd vdd FILL
XFILL_32_CLKBUF1_21 gnd vdd FILL
XFILL_4_INVX1_46 gnd vdd FILL
XFILL_12_NAND3X1_76 gnd vdd FILL
XFILL_32_CLKBUF1_32 gnd vdd FILL
XFILL_12_NAND3X1_87 gnd vdd FILL
XFILL_5_AND2X2_5 gnd vdd FILL
XFILL_4_INVX1_57 gnd vdd FILL
XFILL_12_NAND3X1_98 gnd vdd FILL
XFILL_3_BUFX2_4 gnd vdd FILL
XFILL_4_INVX1_68 gnd vdd FILL
XFILL_13_AOI22X1_7 gnd vdd FILL
XFILL_4_INVX1_79 gnd vdd FILL
XFILL_17_AOI22X1_6 gnd vdd FILL
XFILL_2_BUFX4_11 gnd vdd FILL
XFILL_62_DFFSR_3 gnd vdd FILL
XFILL_2_BUFX4_22 gnd vdd FILL
XFILL_2_BUFX4_33 gnd vdd FILL
XFILL_2_BUFX4_44 gnd vdd FILL
XFILL_19_DFFSR_15 gnd vdd FILL
XFILL_19_DFFSR_26 gnd vdd FILL
XFILL_2_BUFX4_55 gnd vdd FILL
XFILL_19_DFFSR_37 gnd vdd FILL
XFILL_2_BUFX4_66 gnd vdd FILL
XFILL_2_BUFX4_77 gnd vdd FILL
XFILL_19_DFFSR_48 gnd vdd FILL
XFILL_2_BUFX4_88 gnd vdd FILL
XFILL_3_OAI22X1_17 gnd vdd FILL
XFILL_2_BUFX4_99 gnd vdd FILL
XFILL_19_DFFSR_59 gnd vdd FILL
XFILL_3_OAI22X1_28 gnd vdd FILL
XFILL_3_OAI22X1_39 gnd vdd FILL
XFILL_47_5_2 gnd vdd FILL
XFILL_7_OAI21X1_19 gnd vdd FILL
XFILL_59_DFFSR_14 gnd vdd FILL
XFILL_16_AOI22X1_10 gnd vdd FILL
XFILL_59_DFFSR_25 gnd vdd FILL
XFILL_46_0_1 gnd vdd FILL
XFILL_59_DFFSR_36 gnd vdd FILL
XFILL_59_DFFSR_47 gnd vdd FILL
XFILL_59_DFFSR_58 gnd vdd FILL
XFILL_59_DFFSR_69 gnd vdd FILL
XFILL_20_MUX2X1_9 gnd vdd FILL
XFILL_2_NAND3X1_60 gnd vdd FILL
XFILL_2_NAND3X1_71 gnd vdd FILL
XFILL_10_DFFSR_102 gnd vdd FILL
XFILL_2_NAND3X1_82 gnd vdd FILL
XFILL_6_NAND2X1_40 gnd vdd FILL
XFILL_2_NAND3X1_93 gnd vdd FILL
XFILL_6_NAND2X1_51 gnd vdd FILL
XFILL_10_DFFSR_113 gnd vdd FILL
XFILL_10_DFFSR_124 gnd vdd FILL
XFILL_27_DFFSR_6 gnd vdd FILL
XFILL_6_NAND2X1_62 gnd vdd FILL
XFILL_6_NAND2X1_73 gnd vdd FILL
XFILL_10_DFFSR_135 gnd vdd FILL
XFILL_84_DFFSR_7 gnd vdd FILL
XFILL_10_DFFSR_146 gnd vdd FILL
XFILL_28_DFFSR_13 gnd vdd FILL
XFILL_6_NAND2X1_84 gnd vdd FILL
XFILL_10_DFFSR_157 gnd vdd FILL
XFILL_28_DFFSR_24 gnd vdd FILL
XFILL_6_NAND2X1_95 gnd vdd FILL
XFILL_28_DFFSR_35 gnd vdd FILL
XFILL_10_DFFSR_168 gnd vdd FILL
XFILL_28_DFFSR_46 gnd vdd FILL
XFILL_3_INVX2_4 gnd vdd FILL
XFILL_10_DFFSR_179 gnd vdd FILL
XFILL_28_DFFSR_57 gnd vdd FILL
XFILL_14_DFFSR_101 gnd vdd FILL
XFILL_30_4_2 gnd vdd FILL
XFILL_28_DFFSR_68 gnd vdd FILL
XFILL_14_CLKBUF1_15 gnd vdd FILL
XFILL_14_DFFSR_112 gnd vdd FILL
XFILL_28_DFFSR_79 gnd vdd FILL
XFILL_14_CLKBUF1_26 gnd vdd FILL
XFILL_14_DFFSR_123 gnd vdd FILL
XFILL_14_CLKBUF1_37 gnd vdd FILL
XFILL_14_DFFSR_134 gnd vdd FILL
XFILL_68_DFFSR_12 gnd vdd FILL
XFILL_14_DFFSR_145 gnd vdd FILL
XFILL_14_DFFSR_156 gnd vdd FILL
XFILL_68_DFFSR_23 gnd vdd FILL
XFILL_14_DFFSR_167 gnd vdd FILL
XFILL_68_DFFSR_34 gnd vdd FILL
XFILL_14_DFFSR_178 gnd vdd FILL
XFILL_68_DFFSR_45 gnd vdd FILL
XFILL_68_DFFSR_56 gnd vdd FILL
XFILL_68_DFFSR_67 gnd vdd FILL
XFILL_18_DFFSR_100 gnd vdd FILL
XFILL_14_DFFSR_189 gnd vdd FILL
XFILL_18_DFFSR_111 gnd vdd FILL
XFILL_68_DFFSR_78 gnd vdd FILL
XFILL_1_INVX1_2 gnd vdd FILL
XFILL_18_DFFSR_122 gnd vdd FILL
XFILL_68_DFFSR_89 gnd vdd FILL
XFILL_18_DFFSR_133 gnd vdd FILL
XFILL_18_DFFSR_144 gnd vdd FILL
XFILL_18_DFFSR_155 gnd vdd FILL
XCLKBUF1_1 BUFX4_10/Y gnd CLKBUF1_1/Y vdd CLKBUF1
XFILL_18_DFFSR_166 gnd vdd FILL
XFILL_7_CLKBUF1_9 gnd vdd FILL
XFILL_18_DFFSR_177 gnd vdd FILL
XFILL_10_NOR3X1_13 gnd vdd FILL
XFILL_37_DFFSR_11 gnd vdd FILL
XFILL_18_DFFSR_188 gnd vdd FILL
XFILL_10_NOR3X1_24 gnd vdd FILL
XFILL_37_DFFSR_22 gnd vdd FILL
XFILL_10_NOR3X1_35 gnd vdd FILL
XFILL_18_DFFSR_199 gnd vdd FILL
XFILL_10_NOR3X1_46 gnd vdd FILL
XFILL_37_DFFSR_33 gnd vdd FILL
XFILL_60_DFFSR_202 gnd vdd FILL
XFILL_37_DFFSR_44 gnd vdd FILL
XFILL_37_DFFSR_55 gnd vdd FILL
XFILL_60_DFFSR_213 gnd vdd FILL
XFILL_37_DFFSR_66 gnd vdd FILL
XFILL_60_DFFSR_224 gnd vdd FILL
XFILL_37_DFFSR_77 gnd vdd FILL
XFILL_60_DFFSR_235 gnd vdd FILL
XFILL_3_BUFX4_104 gnd vdd FILL
XFILL_60_DFFSR_246 gnd vdd FILL
XFILL_37_DFFSR_88 gnd vdd FILL
XFILL_14_NOR3X1_12 gnd vdd FILL
XFILL_37_DFFSR_99 gnd vdd FILL
XFILL_77_DFFSR_10 gnd vdd FILL
XFILL_60_DFFSR_257 gnd vdd FILL
XFILL_60_DFFSR_268 gnd vdd FILL
XFILL_77_DFFSR_21 gnd vdd FILL
XFILL_14_NOR3X1_23 gnd vdd FILL
XFILL_14_NOR3X1_34 gnd vdd FILL
XFILL_77_DFFSR_32 gnd vdd FILL
XFILL_64_DFFSR_201 gnd vdd FILL
XFILL_14_NOR3X1_45 gnd vdd FILL
XFILL_77_DFFSR_43 gnd vdd FILL
XFILL_64_DFFSR_212 gnd vdd FILL
XFILL_77_DFFSR_54 gnd vdd FILL
XFILL_77_DFFSR_65 gnd vdd FILL
XFILL_64_DFFSR_223 gnd vdd FILL
XFILL_77_DFFSR_76 gnd vdd FILL
XFILL_64_DFFSR_234 gnd vdd FILL
XFILL_38_5_2 gnd vdd FILL
XFILL_7_BUFX4_103 gnd vdd FILL
XFILL_77_DFFSR_87 gnd vdd FILL
XFILL_64_DFFSR_245 gnd vdd FILL
XFILL_18_NOR3X1_11 gnd vdd FILL
XFILL_4_CLKBUF1_10 gnd vdd FILL
XFILL_77_DFFSR_98 gnd vdd FILL
XFILL_37_0_1 gnd vdd FILL
XFILL_64_DFFSR_256 gnd vdd FILL
XFILL_4_CLKBUF1_21 gnd vdd FILL
XFILL_64_DFFSR_267 gnd vdd FILL
XFILL_18_NOR3X1_22 gnd vdd FILL
XFILL_4_CLKBUF1_32 gnd vdd FILL
XFILL_18_NOR3X1_33 gnd vdd FILL
XFILL_0_INVX1_50 gnd vdd FILL
XFILL_68_DFFSR_200 gnd vdd FILL
XFILL_18_NOR3X1_44 gnd vdd FILL
XFILL_0_INVX1_61 gnd vdd FILL
XFILL_68_DFFSR_211 gnd vdd FILL
XFILL_12_MUX2X1_106 gnd vdd FILL
XFILL_0_INVX1_72 gnd vdd FILL
XFILL_12_MUX2X1_117 gnd vdd FILL
XFILL_68_DFFSR_222 gnd vdd FILL
XFILL_0_INVX1_83 gnd vdd FILL
XFILL_46_DFFSR_20 gnd vdd FILL
XFILL_12_MUX2X1_128 gnd vdd FILL
XFILL_0_INVX1_94 gnd vdd FILL
XFILL_68_DFFSR_233 gnd vdd FILL
XFILL_46_DFFSR_31 gnd vdd FILL
XFILL_17_NOR3X1_6 gnd vdd FILL
XFILL_46_DFFSR_42 gnd vdd FILL
XFILL_12_MUX2X1_139 gnd vdd FILL
XFILL_68_DFFSR_244 gnd vdd FILL
XFILL_68_DFFSR_255 gnd vdd FILL
XFILL_46_DFFSR_53 gnd vdd FILL
XFILL_23_CLKBUF1_7 gnd vdd FILL
XFILL_46_DFFSR_64 gnd vdd FILL
XFILL_68_DFFSR_266 gnd vdd FILL
XFILL_46_DFFSR_75 gnd vdd FILL
XFILL_46_DFFSR_86 gnd vdd FILL
XFILL_13_OAI21X1_11 gnd vdd FILL
XFILL_46_DFFSR_97 gnd vdd FILL
XFILL_1_NOR2X1_17 gnd vdd FILL
XFILL_1_NOR2X1_28 gnd vdd FILL
XFILL_13_OAI21X1_22 gnd vdd FILL
XFILL_86_DFFSR_30 gnd vdd FILL
XFILL_1_NOR2X1_39 gnd vdd FILL
XFILL_13_OAI21X1_33 gnd vdd FILL
XFILL_21_4_2 gnd vdd FILL
XFILL_86_DFFSR_41 gnd vdd FILL
XFILL_13_OAI21X1_44 gnd vdd FILL
XFILL_2_NOR2X1_150 gnd vdd FILL
XFILL_86_DFFSR_52 gnd vdd FILL
XFILL_2_NOR2X1_161 gnd vdd FILL
XFILL_86_DFFSR_63 gnd vdd FILL
XFILL_2_NOR2X1_172 gnd vdd FILL
XFILL_27_CLKBUF1_6 gnd vdd FILL
XFILL_86_DFFSR_74 gnd vdd FILL
XFILL_2_NOR2X1_183 gnd vdd FILL
XFILL_15_DFFSR_30 gnd vdd FILL
XFILL_86_DFFSR_85 gnd vdd FILL
XFILL_2_NOR2X1_194 gnd vdd FILL
XFILL_15_DFFSR_41 gnd vdd FILL
XFILL_86_DFFSR_96 gnd vdd FILL
XFILL_15_DFFSR_52 gnd vdd FILL
XFILL_5_NOR2X1_16 gnd vdd FILL
XFILL_5_NOR2X1_27 gnd vdd FILL
XFILL_15_DFFSR_63 gnd vdd FILL
XFILL_5_NOR2X1_38 gnd vdd FILL
XFILL_15_DFFSR_74 gnd vdd FILL
XFILL_15_DFFSR_85 gnd vdd FILL
XFILL_5_NOR2X1_49 gnd vdd FILL
XFILL_15_DFFSR_96 gnd vdd FILL
XFILL_55_DFFSR_40 gnd vdd FILL
XFILL_26_NOR3X1_4 gnd vdd FILL
XFILL_55_DFFSR_51 gnd vdd FILL
XFILL_9_NOR2X1_15 gnd vdd FILL
XFILL_9_NOR2X1_26 gnd vdd FILL
XFILL_55_DFFSR_62 gnd vdd FILL
XFILL_9_NOR2X1_37 gnd vdd FILL
XFILL_55_DFFSR_73 gnd vdd FILL
XFILL_9_NOR2X1_48 gnd vdd FILL
XFILL_55_DFFSR_84 gnd vdd FILL
XFILL_55_DFFSR_95 gnd vdd FILL
XFILL_9_NOR2X1_59 gnd vdd FILL
XFILL_2_MUX2X1_101 gnd vdd FILL
XFILL_2_MUX2X1_112 gnd vdd FILL
XFILL_0_NOR2X1_5 gnd vdd FILL
XFILL_2_MUX2X1_123 gnd vdd FILL
XFILL_2_MUX2X1_134 gnd vdd FILL
XFILL_2_MUX2X1_145 gnd vdd FILL
XFILL_2_MUX2X1_156 gnd vdd FILL
XFILL_2_MUX2X1_167 gnd vdd FILL
XFILL_17_OAI22X1_9 gnd vdd FILL
XFILL_24_DFFSR_50 gnd vdd FILL
XFILL_2_MUX2X1_178 gnd vdd FILL
XFILL_24_DFFSR_61 gnd vdd FILL
XFILL_2_MUX2X1_189 gnd vdd FILL
XFILL_24_DFFSR_72 gnd vdd FILL
XFILL_24_DFFSR_83 gnd vdd FILL
XFILL_29_5_2 gnd vdd FILL
XFILL_4_5_2 gnd vdd FILL
XFILL_24_DFFSR_94 gnd vdd FILL
XFILL_31_DFFSR_201 gnd vdd FILL
XFILL_9_NOR3X1_5 gnd vdd FILL
XFILL_31_DFFSR_212 gnd vdd FILL
XFILL_28_0_1 gnd vdd FILL
XFILL_7_BUFX2_5 gnd vdd FILL
XFILL_3_OAI21X1_50 gnd vdd FILL
XFILL_3_0_1 gnd vdd FILL
XFILL_31_DFFSR_223 gnd vdd FILL
XFILL_31_DFFSR_234 gnd vdd FILL
XFILL_31_DFFSR_245 gnd vdd FILL
XFILL_64_DFFSR_60 gnd vdd FILL
XFILL_31_DFFSR_256 gnd vdd FILL
XFILL_64_DFFSR_71 gnd vdd FILL
XFILL_64_DFFSR_82 gnd vdd FILL
XFILL_31_DFFSR_267 gnd vdd FILL
XFILL_64_DFFSR_93 gnd vdd FILL
XFILL_35_DFFSR_200 gnd vdd FILL
XFILL_35_DFFSR_211 gnd vdd FILL
XFILL_35_DFFSR_222 gnd vdd FILL
XFILL_35_DFFSR_233 gnd vdd FILL
XFILL_35_DFFSR_244 gnd vdd FILL
XFILL_66_DFFSR_4 gnd vdd FILL
XFILL_7_DFFSR_40 gnd vdd FILL
XFILL_35_DFFSR_255 gnd vdd FILL
XFILL_7_DFFSR_51 gnd vdd FILL
XFILL_40_7_0 gnd vdd FILL
XFILL_1_MUX2X1_13 gnd vdd FILL
XFILL_7_DFFSR_62 gnd vdd FILL
XFILL_35_DFFSR_266 gnd vdd FILL
XFILL_7_DFFSR_73 gnd vdd FILL
XFILL_1_MUX2X1_24 gnd vdd FILL
XFILL_62_DFFSR_100 gnd vdd FILL
XFILL_1_MUX2X1_35 gnd vdd FILL
XFILL_12_4_2 gnd vdd FILL
XFILL_7_DFFSR_84 gnd vdd FILL
XFILL_39_DFFSR_210 gnd vdd FILL
XFILL_5_OR2X2_1 gnd vdd FILL
XFILL_62_DFFSR_111 gnd vdd FILL
XINVX8_3 din[3] gnd INVX8_3/Y vdd INVX8
XFILL_7_DFFSR_95 gnd vdd FILL
XFILL_33_DFFSR_70 gnd vdd FILL
XFILL_62_DFFSR_122 gnd vdd FILL
XFILL_1_MUX2X1_46 gnd vdd FILL
XFILL_62_DFFSR_133 gnd vdd FILL
XFILL_39_DFFSR_221 gnd vdd FILL
XFILL_33_DFFSR_81 gnd vdd FILL
XFILL_1_MUX2X1_57 gnd vdd FILL
XFILL_33_DFFSR_92 gnd vdd FILL
XFILL_1_MUX2X1_68 gnd vdd FILL
XFILL_39_DFFSR_232 gnd vdd FILL
XFILL_39_DFFSR_243 gnd vdd FILL
XFILL_1_MUX2X1_79 gnd vdd FILL
XFILL_62_DFFSR_144 gnd vdd FILL
XFILL_62_DFFSR_155 gnd vdd FILL
XFILL_39_DFFSR_254 gnd vdd FILL
XFILL_62_DFFSR_166 gnd vdd FILL
XFILL_39_DFFSR_265 gnd vdd FILL
XFILL_62_DFFSR_177 gnd vdd FILL
XFILL_5_MUX2X1_12 gnd vdd FILL
XFILL_5_MUX2X1_23 gnd vdd FILL
XFILL_5_MUX2X1_34 gnd vdd FILL
XFILL_62_DFFSR_188 gnd vdd FILL
XFILL_5_MUX2X1_45 gnd vdd FILL
XFILL_66_DFFSR_110 gnd vdd FILL
XFILL_62_DFFSR_199 gnd vdd FILL
XFILL_5_NAND3X1_15 gnd vdd FILL
XFILL_66_DFFSR_121 gnd vdd FILL
XFILL_73_DFFSR_80 gnd vdd FILL
XFILL_66_DFFSR_132 gnd vdd FILL
XFILL_5_NAND3X1_26 gnd vdd FILL
XFILL_5_MUX2X1_56 gnd vdd FILL
XFILL_66_DFFSR_143 gnd vdd FILL
XFILL_73_DFFSR_91 gnd vdd FILL
XFILL_5_MUX2X1_67 gnd vdd FILL
XFILL_5_MUX2X1_78 gnd vdd FILL
XFILL_5_NAND3X1_37 gnd vdd FILL
XFILL_66_DFFSR_154 gnd vdd FILL
XFILL_5_NAND3X1_48 gnd vdd FILL
XFILL_5_MUX2X1_89 gnd vdd FILL
XFILL_5_NAND3X1_59 gnd vdd FILL
XFILL_66_DFFSR_165 gnd vdd FILL
XFILL_9_MUX2X1_11 gnd vdd FILL
XFILL_66_DFFSR_176 gnd vdd FILL
XFILL_9_NAND2X1_17 gnd vdd FILL
XFILL_9_MUX2X1_22 gnd vdd FILL
XFILL_9_NAND2X1_28 gnd vdd FILL
XFILL_66_DFFSR_187 gnd vdd FILL
XFILL_9_MUX2X1_33 gnd vdd FILL
XFILL_9_NAND2X1_39 gnd vdd FILL
XFILL_66_DFFSR_198 gnd vdd FILL
XFILL_9_MUX2X1_44 gnd vdd FILL
XFILL_9_MUX2X1_55 gnd vdd FILL
XFILL_9_MUX2X1_66 gnd vdd FILL
XFILL_9_MUX2X1_77 gnd vdd FILL
XFILL_9_MUX2X1_88 gnd vdd FILL
XFILL_9_MUX2X1_99 gnd vdd FILL
XFILL_7_INVX2_5 gnd vdd FILL
XFILL_42_DFFSR_90 gnd vdd FILL
XBUFX4_12 BUFX4_3/Y gnd DFFSR_69/R vdd BUFX4
XFILL_19_MUX2X1_170 gnd vdd FILL
XFILL_10_NOR2X1_90 gnd vdd FILL
XBUFX4_23 BUFX4_51/Y gnd BUFX4_23/Y vdd BUFX4
XFILL_19_MUX2X1_181 gnd vdd FILL
XFILL_19_MUX2X1_192 gnd vdd FILL
XBUFX4_34 BUFX4_62/Y gnd DFFSR_55/R vdd BUFX4
XBUFX4_45 BUFX4_3/Y gnd DFFSR_97/R vdd BUFX4
XBUFX4_56 BUFX4_62/Y gnd DFFSR_96/R vdd BUFX4
XBUFX4_67 INVX8_1/Y gnd BUFX4_67/Y vdd BUFX4
XBUFX4_78 INVX8_2/Y gnd BUFX4_78/Y vdd BUFX4
XFILL_19_0_1 gnd vdd FILL
XBUFX4_89 BUFX4_92/A gnd BUFX4_89/Y vdd BUFX4
XFILL_21_MUX2X1_10 gnd vdd FILL
XFILL_21_MUX2X1_21 gnd vdd FILL
XFILL_5_INVX1_3 gnd vdd FILL
XFILL_21_MUX2X1_32 gnd vdd FILL
XFILL_21_MUX2X1_43 gnd vdd FILL
XFILL_21_MUX2X1_54 gnd vdd FILL
XFILL_62_3_2 gnd vdd FILL
XFILL_21_MUX2X1_65 gnd vdd FILL
XFILL_21_MUX2X1_76 gnd vdd FILL
XFILL_21_MUX2X1_87 gnd vdd FILL
XFILL_21_MUX2X1_98 gnd vdd FILL
XFILL_31_7_0 gnd vdd FILL
XFILL_10_4 gnd vdd FILL
XFILL_24_CLKBUF1_16 gnd vdd FILL
XFILL_24_CLKBUF1_27 gnd vdd FILL
XFILL_24_CLKBUF1_38 gnd vdd FILL
XFILL_33_DFFSR_110 gnd vdd FILL
XFILL_10_NAND2X1_1 gnd vdd FILL
XFILL_33_DFFSR_121 gnd vdd FILL
XFILL_33_DFFSR_132 gnd vdd FILL
XFILL_2_AOI21X1_17 gnd vdd FILL
XFILL_2_AOI21X1_28 gnd vdd FILL
XFILL_33_DFFSR_143 gnd vdd FILL
XFILL_2_AOI21X1_39 gnd vdd FILL
XFILL_33_DFFSR_154 gnd vdd FILL
XFILL_33_DFFSR_165 gnd vdd FILL
XFILL_12_OAI22X1_19 gnd vdd FILL
XFILL_33_DFFSR_176 gnd vdd FILL
XFILL_33_DFFSR_187 gnd vdd FILL
XFILL_33_DFFSR_198 gnd vdd FILL
XFILL_5_NOR2X1_105 gnd vdd FILL
XFILL_37_DFFSR_120 gnd vdd FILL
XFILL_37_DFFSR_131 gnd vdd FILL
XFILL_5_NOR2X1_116 gnd vdd FILL
XFILL_37_DFFSR_142 gnd vdd FILL
XFILL_5_NOR2X1_127 gnd vdd FILL
XFILL_5_NOR2X1_138 gnd vdd FILL
XFILL_37_DFFSR_153 gnd vdd FILL
XFILL_5_NOR2X1_149 gnd vdd FILL
XFILL_37_DFFSR_164 gnd vdd FILL
XFILL_37_DFFSR_175 gnd vdd FILL
XFILL_11_NAND3X1_40 gnd vdd FILL
XFILL_37_DFFSR_186 gnd vdd FILL
XFILL_11_NAND3X1_51 gnd vdd FILL
XFILL_11_NAND3X1_62 gnd vdd FILL
XFILL_37_DFFSR_197 gnd vdd FILL
XFILL_11_NAND3X1_73 gnd vdd FILL
XFILL_11_NAND3X1_84 gnd vdd FILL
XFILL_11_NAND3X1_95 gnd vdd FILL
XFILL_31_CLKBUF1_40 gnd vdd FILL
XFILL_53_3_2 gnd vdd FILL
XFILL_22_MUX2X1_107 gnd vdd FILL
XFILL_83_DFFSR_210 gnd vdd FILL
XFILL_22_MUX2X1_118 gnd vdd FILL
XFILL_10_DFFSR_3 gnd vdd FILL
XFILL_22_MUX2X1_129 gnd vdd FILL
XFILL_83_DFFSR_221 gnd vdd FILL
XFILL_10_AOI21X1_6 gnd vdd FILL
XFILL_83_DFFSR_232 gnd vdd FILL
XFILL_83_DFFSR_243 gnd vdd FILL
XFILL_83_DFFSR_254 gnd vdd FILL
XFILL_22_7_0 gnd vdd FILL
XFILL_83_DFFSR_265 gnd vdd FILL
XFILL_19_DFFSR_109 gnd vdd FILL
XFILL_48_DFFSR_1 gnd vdd FILL
XFILL_1_INVX1_17 gnd vdd FILL
XFILL_1_INVX1_28 gnd vdd FILL
XFILL_87_DFFSR_220 gnd vdd FILL
XFILL_1_INVX1_39 gnd vdd FILL
XFILL_14_AOI21X1_5 gnd vdd FILL
XFILL_2_OAI22X1_14 gnd vdd FILL
XFILL_87_DFFSR_231 gnd vdd FILL
XFILL_87_DFFSR_242 gnd vdd FILL
XFILL_2_OAI22X1_25 gnd vdd FILL
XFILL_87_DFFSR_253 gnd vdd FILL
XFILL_2_OAI22X1_36 gnd vdd FILL
XFILL_2_OAI22X1_47 gnd vdd FILL
XFILL_87_DFFSR_264 gnd vdd FILL
XFILL_87_DFFSR_275 gnd vdd FILL
XFILL_6_OAI21X1_16 gnd vdd FILL
XFILL_6_OAI21X1_27 gnd vdd FILL
XFILL_6_OAI21X1_38 gnd vdd FILL
XFILL_6_OAI21X1_49 gnd vdd FILL
XFILL_3_INVX1_170 gnd vdd FILL
XFILL_3_INVX1_181 gnd vdd FILL
XFILL_3_INVX1_192 gnd vdd FILL
XFILL_87_DFFSR_19 gnd vdd FILL
XFILL_32_DFFSR_7 gnd vdd FILL
XFILL_1_NAND3X1_90 gnd vdd FILL
XFILL_16_DFFSR_19 gnd vdd FILL
XFILL_5_NAND2X1_70 gnd vdd FILL
XFILL_5_NAND2X1_81 gnd vdd FILL
XFILL_5_NAND2X1_92 gnd vdd FILL
XFILL_7_INVX1_180 gnd vdd FILL
XFILL_7_INVX1_191 gnd vdd FILL
XFILL_13_CLKBUF1_12 gnd vdd FILL
XFILL_13_CLKBUF1_23 gnd vdd FILL
XFILL_69_DFFSR_209 gnd vdd FILL
XFILL_13_CLKBUF1_34 gnd vdd FILL
XFILL_56_DFFSR_18 gnd vdd FILL
XFILL_56_DFFSR_29 gnd vdd FILL
XFILL_44_3_2 gnd vdd FILL
XFILL_11_NOR2X1_130 gnd vdd FILL
XFILL_11_NOR2X1_141 gnd vdd FILL
XFILL_25_DFFSR_17 gnd vdd FILL
XFILL_25_DFFSR_28 gnd vdd FILL
XFILL_11_NOR2X1_152 gnd vdd FILL
XFILL_25_DFFSR_39 gnd vdd FILL
XFILL_11_NOR2X1_163 gnd vdd FILL
XFILL_11_NOR2X1_174 gnd vdd FILL
XFILL_50_DFFSR_210 gnd vdd FILL
XFILL_11_NOR2X1_185 gnd vdd FILL
XFILL_13_7_0 gnd vdd FILL
XFILL_50_DFFSR_221 gnd vdd FILL
XFILL_11_NOR2X1_196 gnd vdd FILL
XFILL_50_DFFSR_232 gnd vdd FILL
XFILL_50_DFFSR_243 gnd vdd FILL
XFILL_50_DFFSR_254 gnd vdd FILL
XFILL_65_DFFSR_16 gnd vdd FILL
XFILL_65_DFFSR_27 gnd vdd FILL
XFILL_50_DFFSR_265 gnd vdd FILL
XFILL_9_AOI21X1_70 gnd vdd FILL
XFILL_65_DFFSR_38 gnd vdd FILL
XFILL_9_AOI21X1_81 gnd vdd FILL
XFILL_65_DFFSR_49 gnd vdd FILL
XFILL_19_OAI22X1_50 gnd vdd FILL
XFILL_54_DFFSR_220 gnd vdd FILL
XFILL_54_DFFSR_231 gnd vdd FILL
XFILL_54_DFFSR_242 gnd vdd FILL
XFILL_54_DFFSR_253 gnd vdd FILL
XFILL_54_DFFSR_264 gnd vdd FILL
XFILL_54_DFFSR_275 gnd vdd FILL
XFILL_8_DFFSR_18 gnd vdd FILL
XFILL_8_DFFSR_29 gnd vdd FILL
XFILL_3_CLKBUF1_40 gnd vdd FILL
XFILL_11_MUX2X1_103 gnd vdd FILL
XFILL_34_DFFSR_15 gnd vdd FILL
XFILL_11_MUX2X1_114 gnd vdd FILL
XFILL_81_DFFSR_120 gnd vdd FILL
XFILL_34_DFFSR_26 gnd vdd FILL
XFILL_81_DFFSR_131 gnd vdd FILL
XFILL_11_MUX2X1_125 gnd vdd FILL
XFILL_34_DFFSR_37 gnd vdd FILL
XFILL_58_DFFSR_230 gnd vdd FILL
XFILL_11_MUX2X1_136 gnd vdd FILL
XFILL_81_DFFSR_142 gnd vdd FILL
XFILL_58_DFFSR_241 gnd vdd FILL
XFILL_34_DFFSR_48 gnd vdd FILL
XFILL_81_DFFSR_153 gnd vdd FILL
XFILL_58_DFFSR_252 gnd vdd FILL
XFILL_34_DFFSR_59 gnd vdd FILL
XFILL_11_MUX2X1_147 gnd vdd FILL
XFILL_11_MUX2X1_158 gnd vdd FILL
XFILL_58_DFFSR_263 gnd vdd FILL
XFILL_81_DFFSR_164 gnd vdd FILL
XFILL_81_DFFSR_175 gnd vdd FILL
XFILL_13_CLKBUF1_4 gnd vdd FILL
XFILL_11_MUX2X1_169 gnd vdd FILL
XFILL_1_DFFSR_201 gnd vdd FILL
XFILL_58_DFFSR_274 gnd vdd FILL
XFILL_81_DFFSR_186 gnd vdd FILL
XFILL_81_DFFSR_197 gnd vdd FILL
XFILL_1_DFFSR_212 gnd vdd FILL
XFILL_74_DFFSR_14 gnd vdd FILL
XFILL_1_DFFSR_223 gnd vdd FILL
XFILL_74_DFFSR_25 gnd vdd FILL
XFILL_85_DFFSR_130 gnd vdd FILL
XFILL_1_DFFSR_234 gnd vdd FILL
XFILL_74_DFFSR_36 gnd vdd FILL
XFILL_9_3 gnd vdd FILL
XFILL_12_OAI21X1_30 gnd vdd FILL
XFILL_1_DFFSR_245 gnd vdd FILL
XFILL_85_DFFSR_141 gnd vdd FILL
XFILL_17_MUX2X1_4 gnd vdd FILL
XFILL_12_OAI21X1_41 gnd vdd FILL
XFILL_74_DFFSR_47 gnd vdd FILL
XFILL_85_DFFSR_152 gnd vdd FILL
XFILL_74_DFFSR_58 gnd vdd FILL
XFILL_1_DFFSR_256 gnd vdd FILL
XFILL_1_DFFSR_267 gnd vdd FILL
XFILL_74_DFFSR_69 gnd vdd FILL
XFILL_85_DFFSR_163 gnd vdd FILL
XFILL_85_DFFSR_174 gnd vdd FILL
XFILL_17_CLKBUF1_3 gnd vdd FILL
XFILL_65_5 gnd vdd FILL
XFILL_5_DFFSR_200 gnd vdd FILL
XFILL_1_NOR2X1_180 gnd vdd FILL
XFILL_85_DFFSR_185 gnd vdd FILL
XFILL_5_DFFSR_211 gnd vdd FILL
XFILL_1_NOR2X1_191 gnd vdd FILL
XFILL_85_DFFSR_196 gnd vdd FILL
XFILL_5_DFFSR_222 gnd vdd FILL
XFILL_36_DFFSR_209 gnd vdd FILL
XFILL_5_DFFSR_233 gnd vdd FILL
XFILL_58_4 gnd vdd FILL
XFILL_5_DFFSR_244 gnd vdd FILL
XFILL_5_DFFSR_255 gnd vdd FILL
XFILL_43_DFFSR_13 gnd vdd FILL
XFILL_8_BUFX4_70 gnd vdd FILL
XFILL_43_DFFSR_24 gnd vdd FILL
XFILL_5_DFFSR_266 gnd vdd FILL
XFILL_43_DFFSR_35 gnd vdd FILL
XFILL_8_BUFX4_81 gnd vdd FILL
XFILL_8_BUFX4_92 gnd vdd FILL
XFILL_43_DFFSR_46 gnd vdd FILL
XFILL_63_6_0 gnd vdd FILL
XFILL_9_DFFSR_210 gnd vdd FILL
XFILL_63_DFFSR_109 gnd vdd FILL
XFILL_43_DFFSR_57 gnd vdd FILL
XFILL_35_3_2 gnd vdd FILL
XFILL_43_DFFSR_68 gnd vdd FILL
XFILL_9_DFFSR_221 gnd vdd FILL
XFILL_43_DFFSR_79 gnd vdd FILL
XFILL_9_DFFSR_232 gnd vdd FILL
XFILL_9_DFFSR_243 gnd vdd FILL
XFILL_9_DFFSR_254 gnd vdd FILL
XFILL_83_DFFSR_12 gnd vdd FILL
XFILL_10_NAND3X1_108 gnd vdd FILL
XFILL_9_DFFSR_265 gnd vdd FILL
XFILL_83_DFFSR_23 gnd vdd FILL
XFILL_10_NAND3X1_119 gnd vdd FILL
XFILL_83_DFFSR_34 gnd vdd FILL
XFILL_83_DFFSR_45 gnd vdd FILL
XFILL_83_DFFSR_56 gnd vdd FILL
XFILL_1_MUX2X1_120 gnd vdd FILL
XFILL_67_DFFSR_108 gnd vdd FILL
XFILL_12_DFFSR_12 gnd vdd FILL
XFILL_83_DFFSR_67 gnd vdd FILL
XFILL_67_DFFSR_119 gnd vdd FILL
XFILL_1_MUX2X1_131 gnd vdd FILL
XFILL_12_DFFSR_23 gnd vdd FILL
XFILL_83_DFFSR_78 gnd vdd FILL
XFILL_1_MUX2X1_142 gnd vdd FILL
XFILL_12_DFFSR_34 gnd vdd FILL
XFILL_83_DFFSR_89 gnd vdd FILL
XFILL_1_MUX2X1_153 gnd vdd FILL
XFILL_12_DFFSR_45 gnd vdd FILL
XFILL_12_DFFSR_56 gnd vdd FILL
XFILL_1_MUX2X1_164 gnd vdd FILL
XFILL_14_NAND3X1_17 gnd vdd FILL
XFILL_10_OAI21X1_9 gnd vdd FILL
XFILL_1_MUX2X1_175 gnd vdd FILL
XFILL_12_DFFSR_67 gnd vdd FILL
XFILL_14_NAND3X1_28 gnd vdd FILL
XFILL_12_DFFSR_78 gnd vdd FILL
XFILL_1_MUX2X1_186 gnd vdd FILL
XFILL_14_NAND3X1_39 gnd vdd FILL
XFILL_12_DFFSR_89 gnd vdd FILL
XFILL_52_DFFSR_11 gnd vdd FILL
XFILL_52_DFFSR_22 gnd vdd FILL
XFILL_34_CLKBUF1_17 gnd vdd FILL
XFILL_34_CLKBUF1_28 gnd vdd FILL
XFILL_11_NOR2X1_11 gnd vdd FILL
XFILL_52_DFFSR_33 gnd vdd FILL
XFILL_23_NOR3X1_8 gnd vdd FILL
XFILL_21_DFFSR_220 gnd vdd FILL
XFILL_11_NOR2X1_22 gnd vdd FILL
XFILL_52_DFFSR_44 gnd vdd FILL
XFILL_34_CLKBUF1_39 gnd vdd FILL
XFILL_52_DFFSR_55 gnd vdd FILL
XFILL_2_AOI22X1_5 gnd vdd FILL
XFILL_11_NOR2X1_33 gnd vdd FILL
XFILL_21_DFFSR_231 gnd vdd FILL
XFILL_21_DFFSR_242 gnd vdd FILL
XFILL_11_NOR2X1_44 gnd vdd FILL
XFILL_14_OAI21X1_8 gnd vdd FILL
XFILL_52_DFFSR_66 gnd vdd FILL
XFILL_21_DFFSR_253 gnd vdd FILL
XFILL_52_DFFSR_77 gnd vdd FILL
XFILL_11_NOR2X1_55 gnd vdd FILL
XFILL_11_NOR2X1_66 gnd vdd FILL
XFILL_52_DFFSR_88 gnd vdd FILL
XFILL_21_DFFSR_264 gnd vdd FILL
XFILL_21_DFFSR_275 gnd vdd FILL
XFILL_11_NOR2X1_77 gnd vdd FILL
XFILL_52_DFFSR_99 gnd vdd FILL
XFILL_2_INVX1_204 gnd vdd FILL
XFILL_11_NOR2X1_88 gnd vdd FILL
XFILL_2_INVX1_215 gnd vdd FILL
XFILL_1_DFFSR_6 gnd vdd FILL
XFILL_9_MUX2X1_3 gnd vdd FILL
XFILL_11_NOR2X1_99 gnd vdd FILL
XFILL_2_INVX1_226 gnd vdd FILL
XFILL_14_DFFSR_4 gnd vdd FILL
XFILL_6_AOI22X1_4 gnd vdd FILL
XFILL_25_DFFSR_230 gnd vdd FILL
XFILL_21_DFFSR_10 gnd vdd FILL
XFILL_21_DFFSR_21 gnd vdd FILL
XFILL_25_DFFSR_241 gnd vdd FILL
XFILL_71_DFFSR_5 gnd vdd FILL
XFILL_25_DFFSR_252 gnd vdd FILL
XFILL_21_DFFSR_32 gnd vdd FILL
XFILL_25_DFFSR_263 gnd vdd FILL
XFILL_21_DFFSR_43 gnd vdd FILL
XFILL_25_DFFSR_274 gnd vdd FILL
XFILL_6_INVX1_203 gnd vdd FILL
XFILL_21_DFFSR_54 gnd vdd FILL
XFILL_22_MUX2X1_19 gnd vdd FILL
XFILL_21_DFFSR_65 gnd vdd FILL
XFILL_21_DFFSR_76 gnd vdd FILL
XFILL_6_INVX1_214 gnd vdd FILL
XFILL_6_INVX1_225 gnd vdd FILL
XFILL_52_DFFSR_130 gnd vdd FILL
XFILL_21_DFFSR_87 gnd vdd FILL
XFILL_21_DFFSR_98 gnd vdd FILL
XFILL_52_DFFSR_141 gnd vdd FILL
XFILL_6_NOR3X1_9 gnd vdd FILL
XFILL_61_DFFSR_20 gnd vdd FILL
XFILL_29_DFFSR_240 gnd vdd FILL
XFILL_52_DFFSR_152 gnd vdd FILL
XFILL_29_DFFSR_251 gnd vdd FILL
XFILL_61_DFFSR_31 gnd vdd FILL
XFILL_29_DFFSR_262 gnd vdd FILL
XFILL_52_DFFSR_163 gnd vdd FILL
XFILL_52_DFFSR_174 gnd vdd FILL
XFILL_61_DFFSR_42 gnd vdd FILL
XFILL_61_DFFSR_53 gnd vdd FILL
XFILL_29_DFFSR_273 gnd vdd FILL
XFILL_52_DFFSR_185 gnd vdd FILL
XFILL_61_DFFSR_64 gnd vdd FILL
XFILL_61_DFFSR_75 gnd vdd FILL
XFILL_52_DFFSR_196 gnd vdd FILL
XFILL_61_DFFSR_86 gnd vdd FILL
XFILL_4_NAND3X1_12 gnd vdd FILL
XFILL_4_NAND3X1_23 gnd vdd FILL
XFILL_56_DFFSR_140 gnd vdd FILL
XFILL_4_NAND3X1_34 gnd vdd FILL
XFILL_61_DFFSR_97 gnd vdd FILL
XFILL_54_6_0 gnd vdd FILL
XFILL_56_DFFSR_151 gnd vdd FILL
XFILL_4_DFFSR_11 gnd vdd FILL
XFILL_4_NAND3X1_45 gnd vdd FILL
XFILL_26_3_2 gnd vdd FILL
XFILL_56_DFFSR_162 gnd vdd FILL
XFILL_8_NAND2X1_14 gnd vdd FILL
XFILL_4_DFFSR_22 gnd vdd FILL
XFILL_1_3_2 gnd vdd FILL
XFILL_4_NAND3X1_56 gnd vdd FILL
XFILL_56_DFFSR_173 gnd vdd FILL
XFILL_4_NAND3X1_67 gnd vdd FILL
XFILL_56_DFFSR_184 gnd vdd FILL
XFILL_4_NAND3X1_78 gnd vdd FILL
XFILL_4_DFFSR_33 gnd vdd FILL
XFILL_8_NAND2X1_25 gnd vdd FILL
XFILL_36_DFFSR_8 gnd vdd FILL
XFILL_56_DFFSR_195 gnd vdd FILL
XFILL_8_NAND2X1_36 gnd vdd FILL
XFILL_4_DFFSR_44 gnd vdd FILL
XFILL_30_DFFSR_109 gnd vdd FILL
XFILL_4_DFFSR_55 gnd vdd FILL
XFILL_4_NAND3X1_89 gnd vdd FILL
XFILL_30_DFFSR_30 gnd vdd FILL
XFILL_8_NAND2X1_47 gnd vdd FILL
XFILL_8_NAND2X1_58 gnd vdd FILL
XFILL_4_DFFSR_66 gnd vdd FILL
XFILL_30_DFFSR_41 gnd vdd FILL
XFILL_4_DFFSR_77 gnd vdd FILL
XFILL_8_NAND2X1_69 gnd vdd FILL
XFILL_30_DFFSR_52 gnd vdd FILL
XFILL_30_DFFSR_63 gnd vdd FILL
XFILL_4_DFFSR_88 gnd vdd FILL
XFILL_4_DFFSR_99 gnd vdd FILL
XFILL_30_DFFSR_74 gnd vdd FILL
XFILL_30_DFFSR_85 gnd vdd FILL
XFILL_30_DFFSR_96 gnd vdd FILL
XFILL_3_DFFSR_110 gnd vdd FILL
XFILL_34_DFFSR_108 gnd vdd FILL
XFILL_3_DFFSR_121 gnd vdd FILL
XFILL_70_DFFSR_40 gnd vdd FILL
XFILL_3_DFFSR_132 gnd vdd FILL
XFILL_34_DFFSR_119 gnd vdd FILL
XFILL_70_DFFSR_51 gnd vdd FILL
XFILL_3_DFFSR_143 gnd vdd FILL
XFILL_3_DFFSR_154 gnd vdd FILL
XFILL_70_DFFSR_62 gnd vdd FILL
XFILL_11_AOI21X1_19 gnd vdd FILL
XFILL_3_DFFSR_165 gnd vdd FILL
XFILL_70_DFFSR_73 gnd vdd FILL
XFILL_70_DFFSR_84 gnd vdd FILL
XFILL_3_DFFSR_176 gnd vdd FILL
XFILL_70_DFFSR_95 gnd vdd FILL
XFILL_3_DFFSR_187 gnd vdd FILL
XFILL_3_DFFSR_198 gnd vdd FILL
XFILL_38_DFFSR_107 gnd vdd FILL
XFILL_7_DFFSR_120 gnd vdd FILL
XFILL_7_DFFSR_131 gnd vdd FILL
XFILL_38_DFFSR_118 gnd vdd FILL
XFILL_7_DFFSR_142 gnd vdd FILL
XFILL_11_MUX2X1_40 gnd vdd FILL
XFILL_38_DFFSR_129 gnd vdd FILL
XFILL_7_DFFSR_153 gnd vdd FILL
XFILL_11_MUX2X1_51 gnd vdd FILL
XFILL_11_MUX2X1_62 gnd vdd FILL
XFILL_7_DFFSR_164 gnd vdd FILL
XFILL_11_MUX2X1_73 gnd vdd FILL
XFILL_7_DFFSR_175 gnd vdd FILL
XFILL_10_NOR3X1_3 gnd vdd FILL
XFILL_11_MUX2X1_84 gnd vdd FILL
XFILL_7_DFFSR_186 gnd vdd FILL
XFILL_7_DFFSR_197 gnd vdd FILL
XFILL_11_MUX2X1_95 gnd vdd FILL
XFILL_9_4_2 gnd vdd FILL
XFILL_80_DFFSR_209 gnd vdd FILL
XFILL_15_MUX2X1_50 gnd vdd FILL
XFILL_15_MUX2X1_61 gnd vdd FILL
XFILL_3_NOR3X1_10 gnd vdd FILL
XFILL_15_MUX2X1_72 gnd vdd FILL
XFILL_15_MUX2X1_83 gnd vdd FILL
XFILL_3_NOR3X1_21 gnd vdd FILL
XFILL_15_MUX2X1_94 gnd vdd FILL
XFILL_3_NOR3X1_32 gnd vdd FILL
XFILL_3_NOR3X1_43 gnd vdd FILL
XFILL_23_CLKBUF1_13 gnd vdd FILL
XFILL_84_DFFSR_208 gnd vdd FILL
XFILL_23_CLKBUF1_24 gnd vdd FILL
XFILL_23_CLKBUF1_35 gnd vdd FILL
XFILL_84_DFFSR_219 gnd vdd FILL
XFILL_19_MUX2X1_60 gnd vdd FILL
XFILL_19_MUX2X1_71 gnd vdd FILL
XFILL_19_MUX2X1_82 gnd vdd FILL
XFILL_7_NOR3X1_20 gnd vdd FILL
XFILL_19_MUX2X1_93 gnd vdd FILL
XFILL_7_NOR3X1_31 gnd vdd FILL
XFILL_6_CLKBUF1_17 gnd vdd FILL
XFILL_0_INVX1_103 gnd vdd FILL
XFILL_6_CLKBUF1_28 gnd vdd FILL
XFILL_0_INVX1_114 gnd vdd FILL
XFILL_45_6_0 gnd vdd FILL
XFILL_7_NOR3X1_42 gnd vdd FILL
XFILL_0_INVX1_125 gnd vdd FILL
XFILL_17_3_2 gnd vdd FILL
XFILL_6_CLKBUF1_39 gnd vdd FILL
XFILL_0_INVX1_136 gnd vdd FILL
XFILL_1_AOI21X1_14 gnd vdd FILL
XFILL_0_INVX1_147 gnd vdd FILL
XFILL_23_DFFSR_140 gnd vdd FILL
XFILL_1_AOI21X1_25 gnd vdd FILL
XFILL_1_AOI21X1_36 gnd vdd FILL
XFILL_0_INVX1_158 gnd vdd FILL
XFILL_0_INVX1_169 gnd vdd FILL
XFILL_23_DFFSR_151 gnd vdd FILL
XFILL_1_AOI21X1_47 gnd vdd FILL
XFILL_23_DFFSR_162 gnd vdd FILL
XFILL_1_AOI21X1_58 gnd vdd FILL
XFILL_23_DFFSR_173 gnd vdd FILL
XFILL_11_OAI22X1_16 gnd vdd FILL
XFILL_23_DFFSR_184 gnd vdd FILL
XFILL_4_INVX1_102 gnd vdd FILL
XFILL_1_AOI21X1_69 gnd vdd FILL
XFILL_11_OAI22X1_27 gnd vdd FILL
XFILL_11_OAI22X1_38 gnd vdd FILL
XFILL_4_INVX1_113 gnd vdd FILL
XFILL_23_DFFSR_195 gnd vdd FILL
XFILL_4_INVX1_124 gnd vdd FILL
XFILL_4_NOR2X1_102 gnd vdd FILL
XFILL_4_INVX1_135 gnd vdd FILL
XFILL_11_OAI22X1_49 gnd vdd FILL
XFILL_4_NOR2X1_113 gnd vdd FILL
XFILL_15_OAI21X1_18 gnd vdd FILL
XFILL_4_INVX1_146 gnd vdd FILL
XFILL_4_NOR2X1_124 gnd vdd FILL
XFILL_15_OAI21X1_29 gnd vdd FILL
XFILL_4_INVX1_157 gnd vdd FILL
XFILL_27_DFFSR_150 gnd vdd FILL
XFILL_4_NOR2X1_135 gnd vdd FILL
XFILL_4_NOR2X1_146 gnd vdd FILL
XFILL_4_INVX1_168 gnd vdd FILL
XFILL_27_DFFSR_161 gnd vdd FILL
XFILL_4_INVX1_179 gnd vdd FILL
XFILL_4_NOR2X1_157 gnd vdd FILL
XFILL_27_DFFSR_172 gnd vdd FILL
XFILL_27_DFFSR_183 gnd vdd FILL
XFILL_4_NOR2X1_168 gnd vdd FILL
XFILL_4_NOR2X1_179 gnd vdd FILL
XFILL_27_DFFSR_194 gnd vdd FILL
XFILL_10_NAND3X1_70 gnd vdd FILL
XFILL_11_INVX8_2 gnd vdd FILL
XFILL_2_NOR3X1_2 gnd vdd FILL
XFILL_10_NAND3X1_81 gnd vdd FILL
XFILL_10_NAND3X1_92 gnd vdd FILL
XFILL_23_NOR3X1_40 gnd vdd FILL
XFILL_23_NOR3X1_51 gnd vdd FILL
XFILL_21_MUX2X1_104 gnd vdd FILL
XFILL_21_MUX2X1_115 gnd vdd FILL
XFILL_21_MUX2X1_126 gnd vdd FILL
XFILL_2_OAI22X1_8 gnd vdd FILL
XFILL_21_MUX2X1_137 gnd vdd FILL
XFILL_21_MUX2X1_148 gnd vdd FILL
XFILL_73_DFFSR_240 gnd vdd FILL
XFILL_73_DFFSR_251 gnd vdd FILL
XFILL_21_MUX2X1_159 gnd vdd FILL
XFILL_73_DFFSR_262 gnd vdd FILL
XFILL_53_DFFSR_2 gnd vdd FILL
XFILL_4_MUX2X1_108 gnd vdd FILL
XFILL_0_DFFSR_70 gnd vdd FILL
XFILL_73_DFFSR_273 gnd vdd FILL
XFILL_4_MUX2X1_119 gnd vdd FILL
XFILL_0_DFFSR_81 gnd vdd FILL
XFILL_27_NOR3X1_50 gnd vdd FILL
XFILL_0_DFFSR_92 gnd vdd FILL
XFILL_9_NOR2X1_202 gnd vdd FILL
XFILL_6_OAI22X1_7 gnd vdd FILL
XFILL_1_OAI22X1_11 gnd vdd FILL
XFILL_1_OAI22X1_22 gnd vdd FILL
XFILL_63_2 gnd vdd FILL
XFILL_1_OAI22X1_33 gnd vdd FILL
XFILL_77_DFFSR_250 gnd vdd FILL
XFILL_1_OAI22X1_44 gnd vdd FILL
XFILL_77_DFFSR_261 gnd vdd FILL
XFILL_77_DFFSR_272 gnd vdd FILL
XFILL_32_CLKBUF1_2 gnd vdd FILL
XFILL_5_OAI21X1_13 gnd vdd FILL
XFILL_56_1 gnd vdd FILL
XFILL_5_OAI21X1_24 gnd vdd FILL
XFILL_5_OAI21X1_35 gnd vdd FILL
XFILL_51_DFFSR_208 gnd vdd FILL
XFILL_51_DFFSR_219 gnd vdd FILL
XFILL_5_OAI21X1_46 gnd vdd FILL
XFILL_36_6_0 gnd vdd FILL
XFILL_5_DFFSR_7 gnd vdd FILL
XFILL_55_DFFSR_207 gnd vdd FILL
XFILL_18_DFFSR_5 gnd vdd FILL
XFILL_55_DFFSR_218 gnd vdd FILL
XFILL_55_DFFSR_229 gnd vdd FILL
XFILL_75_DFFSR_6 gnd vdd FILL
XFILL_50_1_2 gnd vdd FILL
XFILL_9_BUFX4_15 gnd vdd FILL
XFILL_11_NAND3X1_109 gnd vdd FILL
XFILL_9_BUFX4_26 gnd vdd FILL
XFILL_9_BUFX4_37 gnd vdd FILL
XFILL_9_BUFX4_48 gnd vdd FILL
XFILL_59_DFFSR_206 gnd vdd FILL
XFILL_82_DFFSR_107 gnd vdd FILL
XFILL_12_CLKBUF1_20 gnd vdd FILL
XFILL_9_BUFX4_59 gnd vdd FILL
XFILL_59_DFFSR_217 gnd vdd FILL
XFILL_12_CLKBUF1_31 gnd vdd FILL
XFILL_82_DFFSR_118 gnd vdd FILL
XFILL_12_CLKBUF1_42 gnd vdd FILL
XFILL_82_DFFSR_129 gnd vdd FILL
XFILL_59_DFFSR_228 gnd vdd FILL
XFILL_59_DFFSR_239 gnd vdd FILL
XFILL_86_DFFSR_106 gnd vdd FILL
XFILL_86_DFFSR_117 gnd vdd FILL
XFILL_86_DFFSR_128 gnd vdd FILL
XFILL_86_DFFSR_139 gnd vdd FILL
XFILL_10_NOR2X1_160 gnd vdd FILL
XFILL_6_DFFSR_209 gnd vdd FILL
XFILL_10_NOR2X1_171 gnd vdd FILL
XFILL_3_NAND3X1_9 gnd vdd FILL
XFILL_10_NOR2X1_182 gnd vdd FILL
XFILL_10_NOR2X1_193 gnd vdd FILL
XFILL_40_DFFSR_240 gnd vdd FILL
XFILL_40_DFFSR_251 gnd vdd FILL
XFILL_40_DFFSR_262 gnd vdd FILL
XFILL_40_DFFSR_273 gnd vdd FILL
XFILL_7_NAND3X1_8 gnd vdd FILL
XFILL_58_2_2 gnd vdd FILL
XFILL_44_DFFSR_250 gnd vdd FILL
XFILL_44_DFFSR_261 gnd vdd FILL
XFILL_13_BUFX4_20 gnd vdd FILL
XFILL_13_BUFX4_31 gnd vdd FILL
XFILL_44_DFFSR_272 gnd vdd FILL
XFILL_13_BUFX4_42 gnd vdd FILL
XFILL_27_6_0 gnd vdd FILL
XFILL_12_BUFX4_5 gnd vdd FILL
XFILL_10_MUX2X1_100 gnd vdd FILL
XFILL_2_6_0 gnd vdd FILL
XFILL_10_MUX2X1_111 gnd vdd FILL
XFILL_13_BUFX4_53 gnd vdd FILL
XFILL_10_MUX2X1_122 gnd vdd FILL
XFILL_13_BUFX4_64 gnd vdd FILL
XFILL_10_MUX2X1_133 gnd vdd FILL
XFILL_13_BUFX4_75 gnd vdd FILL
XFILL_10_MUX2X1_144 gnd vdd FILL
XFILL_13_BUFX4_86 gnd vdd FILL
XFILL_13_BUFX4_97 gnd vdd FILL
XFILL_71_DFFSR_150 gnd vdd FILL
XFILL_71_DFFSR_161 gnd vdd FILL
XFILL_10_MUX2X1_155 gnd vdd FILL
XFILL_48_DFFSR_260 gnd vdd FILL
XFILL_48_DFFSR_271 gnd vdd FILL
XFILL_71_DFFSR_172 gnd vdd FILL
XFILL_10_MUX2X1_166 gnd vdd FILL
XFILL_71_DFFSR_183 gnd vdd FILL
XFILL_10_MUX2X1_177 gnd vdd FILL
XFILL_10_MUX2X1_188 gnd vdd FILL
XFILL_71_DFFSR_194 gnd vdd FILL
XFILL_22_DFFSR_207 gnd vdd FILL
XFILL_41_1_2 gnd vdd FILL
XFILL_22_DFFSR_218 gnd vdd FILL
XFILL_22_DFFSR_229 gnd vdd FILL
XFILL_75_DFFSR_160 gnd vdd FILL
XFILL_75_DFFSR_171 gnd vdd FILL
XFILL_75_DFFSR_182 gnd vdd FILL
XFILL_75_DFFSR_193 gnd vdd FILL
XFILL_10_5_0 gnd vdd FILL
XFILL_26_DFFSR_206 gnd vdd FILL
XAOI22X1_5 INVX1_120/Y NOR2X1_18/A NOR2X1_15/A INVX1_121/Y gnd AOI22X1_5/Y vdd AOI22X1
XFILL_26_DFFSR_217 gnd vdd FILL
XFILL_26_DFFSR_228 gnd vdd FILL
XFILL_31_DFFSR_19 gnd vdd FILL
XFILL_26_DFFSR_239 gnd vdd FILL
XFILL_7_INVX1_10 gnd vdd FILL
XFILL_7_INVX1_21 gnd vdd FILL
XFILL_79_DFFSR_170 gnd vdd FILL
XFILL_7_INVX1_32 gnd vdd FILL
XINVX1_204 DFFSR_88/Q gnd INVX1_204/Y vdd INVX1
XINVX1_215 DFFSR_67/Q gnd INVX1_215/Y vdd INVX1
XFILL_7_INVX1_43 gnd vdd FILL
XFILL_8_AND2X2_2 gnd vdd FILL
XFILL_79_DFFSR_181 gnd vdd FILL
XFILL_7_INVX1_54 gnd vdd FILL
XFILL_79_DFFSR_192 gnd vdd FILL
XINVX1_226 DFFSR_61/Q gnd INVX1_226/Y vdd INVX1
XFILL_53_DFFSR_106 gnd vdd FILL
XFILL_7_INVX1_65 gnd vdd FILL
XFILL_53_DFFSR_117 gnd vdd FILL
XFILL_7_INVX1_76 gnd vdd FILL
XFILL_53_DFFSR_128 gnd vdd FILL
XFILL_7_INVX1_87 gnd vdd FILL
XFILL_53_DFFSR_139 gnd vdd FILL
XFILL_7_INVX1_98 gnd vdd FILL
XFILL_71_DFFSR_18 gnd vdd FILL
XFILL_71_DFFSR_29 gnd vdd FILL
XFILL_14_MUX2X1_8 gnd vdd FILL
XFILL_57_DFFSR_105 gnd vdd FILL
XFILL_57_DFFSR_116 gnd vdd FILL
XFILL_57_DFFSR_127 gnd vdd FILL
XFILL_57_DFFSR_138 gnd vdd FILL
XFILL_0_MUX2X1_150 gnd vdd FILL
XFILL_0_MUX2X1_161 gnd vdd FILL
XFILL_57_DFFSR_149 gnd vdd FILL
XFILL_13_NAND3X1_14 gnd vdd FILL
XFILL_5_BUFX4_30 gnd vdd FILL
XFILL_0_MUX2X1_172 gnd vdd FILL
XNAND2X1_15 INVX2_1/A INVX1_8/A gnd MUX2X1_99/S vdd NAND2X1
XFILL_5_BUFX4_41 gnd vdd FILL
XFILL_49_2_2 gnd vdd FILL
XFILL_13_NAND3X1_25 gnd vdd FILL
XNAND2X1_26 AND2X2_6/B AND2X2_6/A gnd NOR2X1_41/B vdd NAND2X1
XFILL_5_BUFX4_52 gnd vdd FILL
XFILL_13_NAND3X1_36 gnd vdd FILL
XNAND2X1_37 BUFX4_89/Y AND2X2_3/Y gnd OAI22X1_50/D vdd NAND2X1
XFILL_0_MUX2X1_183 gnd vdd FILL
XFILL_5_BUFX4_63 gnd vdd FILL
XNAND2X1_48 BUFX4_7/Y NOR2X1_44/Y gnd NOR2X1_51/B vdd NAND2X1
XFILL_0_MUX2X1_194 gnd vdd FILL
XFILL_13_NAND3X1_47 gnd vdd FILL
XFILL_0_DFFSR_109 gnd vdd FILL
XFILL_13_NAND3X1_58 gnd vdd FILL
XNAND2X1_59 BUFX4_104/Y NOR2X1_30/Y gnd OAI21X1_7/B vdd NAND2X1
XFILL_40_DFFSR_17 gnd vdd FILL
XFILL_13_NAND3X1_69 gnd vdd FILL
XFILL_40_DFFSR_28 gnd vdd FILL
XFILL_5_BUFX4_74 gnd vdd FILL
XFILL_15_INVX8_3 gnd vdd FILL
XFILL_5_BUFX4_85 gnd vdd FILL
XFILL_40_DFFSR_39 gnd vdd FILL
XFILL_33_CLKBUF1_14 gnd vdd FILL
XFILL_33_CLKBUF1_25 gnd vdd FILL
XFILL_5_BUFX4_96 gnd vdd FILL
XFILL_33_CLKBUF1_36 gnd vdd FILL
XFILL_18_6_0 gnd vdd FILL
XFILL_11_DFFSR_250 gnd vdd FILL
XFILL_11_DFFSR_261 gnd vdd FILL
XFILL_4_DFFSR_108 gnd vdd FILL
XFILL_11_DFFSR_272 gnd vdd FILL
XFILL_80_DFFSR_16 gnd vdd FILL
XFILL_80_DFFSR_27 gnd vdd FILL
XFILL_4_DFFSR_119 gnd vdd FILL
XFILL_80_DFFSR_38 gnd vdd FILL
XFILL_80_DFFSR_49 gnd vdd FILL
XFILL_23_MUX2X1_6 gnd vdd FILL
XFILL_60_4_0 gnd vdd FILL
XFILL_28_5 gnd vdd FILL
XFILL_15_DFFSR_260 gnd vdd FILL
XFILL_32_1_2 gnd vdd FILL
XFILL_57_DFFSR_3 gnd vdd FILL
XFILL_15_DFFSR_271 gnd vdd FILL
XFILL_8_DFFSR_107 gnd vdd FILL
XFILL_7_NOR2X1_9 gnd vdd FILL
XFILL_12_MUX2X1_16 gnd vdd FILL
XFILL_8_DFFSR_118 gnd vdd FILL
XFILL_8_DFFSR_129 gnd vdd FILL
XFILL_12_MUX2X1_27 gnd vdd FILL
XFILL_12_MUX2X1_38 gnd vdd FILL
XFILL_3_AOI21X1_3 gnd vdd FILL
XFILL_12_MUX2X1_49 gnd vdd FILL
XFILL_42_DFFSR_160 gnd vdd FILL
XFILL_19_DFFSR_270 gnd vdd FILL
XFILL_42_DFFSR_171 gnd vdd FILL
XFILL_42_DFFSR_182 gnd vdd FILL
XFILL_42_DFFSR_193 gnd vdd FILL
XFILL_16_MUX2X1_15 gnd vdd FILL
XFILL_16_MUX2X1_26 gnd vdd FILL
XFILL_16_MUX2X1_37 gnd vdd FILL
XFILL_3_NAND3X1_20 gnd vdd FILL
XFILL_7_AOI21X1_2 gnd vdd FILL
XFILL_16_MUX2X1_48 gnd vdd FILL
XFILL_3_NAND3X1_31 gnd vdd FILL
XFILL_16_MUX2X1_59 gnd vdd FILL
XFILL_3_NAND3X1_42 gnd vdd FILL
XFILL_6_MUX2X1_7 gnd vdd FILL
XNOR3X1_3 NOR3X1_3/A NOR3X1_3/B NOR3X1_3/C gnd NOR3X1_3/Y vdd NOR3X1
XFILL_7_NAND2X1_11 gnd vdd FILL
XFILL_3_NAND3X1_53 gnd vdd FILL
XFILL_4_NOR3X1_19 gnd vdd FILL
XFILL_46_DFFSR_170 gnd vdd FILL
XFILL_3_NAND3X1_64 gnd vdd FILL
XFILL_3_NAND3X1_75 gnd vdd FILL
XFILL_7_NAND2X1_22 gnd vdd FILL
XFILL_46_DFFSR_181 gnd vdd FILL
XFILL_41_DFFSR_9 gnd vdd FILL
XFILL_3_NAND3X1_86 gnd vdd FILL
XFILL_46_DFFSR_192 gnd vdd FILL
XFILL_7_NAND2X1_33 gnd vdd FILL
XFILL_20_DFFSR_106 gnd vdd FILL
XFILL_9_DFFSR_8 gnd vdd FILL
XFILL_7_NAND2X1_44 gnd vdd FILL
XFILL_7_NAND2X1_55 gnd vdd FILL
XFILL_3_NAND3X1_97 gnd vdd FILL
XFILL_20_DFFSR_117 gnd vdd FILL
XFILL_7_NAND2X1_66 gnd vdd FILL
XFILL_20_DFFSR_128 gnd vdd FILL
XFILL_20_DFFSR_139 gnd vdd FILL
XFILL_7_NAND2X1_77 gnd vdd FILL
XFILL_79_DFFSR_7 gnd vdd FILL
XFILL_7_NAND2X1_88 gnd vdd FILL
XFILL_8_NOR3X1_18 gnd vdd FILL
XFILL_8_NOR3X1_29 gnd vdd FILL
XFILL_24_DFFSR_105 gnd vdd FILL
XFILL_15_CLKBUF1_19 gnd vdd FILL
XFILL_24_DFFSR_116 gnd vdd FILL
XFILL_24_DFFSR_127 gnd vdd FILL
XFILL_24_DFFSR_138 gnd vdd FILL
XFILL_24_DFFSR_149 gnd vdd FILL
XFILL_10_AOI21X1_16 gnd vdd FILL
XFILL_10_AOI21X1_27 gnd vdd FILL
XFILL_10_AOI21X1_38 gnd vdd FILL
XFILL_10_AOI21X1_49 gnd vdd FILL
XFILL_28_DFFSR_104 gnd vdd FILL
XFILL_1_DFFSR_15 gnd vdd FILL
XFILL_1_DFFSR_26 gnd vdd FILL
XFILL_11_NOR2X1_3 gnd vdd FILL
XFILL_28_DFFSR_115 gnd vdd FILL
XFILL_1_DFFSR_37 gnd vdd FILL
XFILL_28_DFFSR_126 gnd vdd FILL
XFILL_28_DFFSR_137 gnd vdd FILL
XFILL_1_DFFSR_48 gnd vdd FILL
XFILL_28_DFFSR_148 gnd vdd FILL
XFILL_1_DFFSR_59 gnd vdd FILL
XFILL_28_DFFSR_159 gnd vdd FILL
XFILL_20_NOR3X1_17 gnd vdd FILL
XFILL_3_INVX1_80 gnd vdd FILL
XFILL_20_NOR3X1_28 gnd vdd FILL
XFILL_3_INVX1_91 gnd vdd FILL
XFILL_51_4_0 gnd vdd FILL
XFILL_20_NOR3X1_39 gnd vdd FILL
XFILL_70_DFFSR_206 gnd vdd FILL
XFILL_23_1_2 gnd vdd FILL
XFILL_70_DFFSR_217 gnd vdd FILL
XFILL_49_DFFSR_50 gnd vdd FILL
XFILL_70_DFFSR_228 gnd vdd FILL
XFILL_49_DFFSR_61 gnd vdd FILL
XFILL_10_MUX2X1_1 gnd vdd FILL
XFILL_70_DFFSR_239 gnd vdd FILL
XFILL_49_DFFSR_72 gnd vdd FILL
XFILL_49_DFFSR_83 gnd vdd FILL
XFILL_24_NOR3X1_16 gnd vdd FILL
XFILL_49_DFFSR_94 gnd vdd FILL
XFILL_24_NOR3X1_27 gnd vdd FILL
XFILL_24_NOR3X1_38 gnd vdd FILL
XFILL_22_CLKBUF1_10 gnd vdd FILL
XFILL_22_CLKBUF1_21 gnd vdd FILL
XFILL_24_NOR3X1_49 gnd vdd FILL
XFILL_74_DFFSR_205 gnd vdd FILL
XFILL_22_CLKBUF1_32 gnd vdd FILL
XFILL_74_DFFSR_216 gnd vdd FILL
XFILL_74_DFFSR_227 gnd vdd FILL
XFILL_74_DFFSR_238 gnd vdd FILL
XFILL_74_DFFSR_249 gnd vdd FILL
XFILL_28_NOR3X1_15 gnd vdd FILL
XFILL_3_BUFX4_8 gnd vdd FILL
XFILL_5_CLKBUF1_14 gnd vdd FILL
XFILL_5_CLKBUF1_25 gnd vdd FILL
XFILL_28_NOR3X1_26 gnd vdd FILL
XFILL_18_DFFSR_60 gnd vdd FILL
XFILL_5_CLKBUF1_36 gnd vdd FILL
XFILL_18_DFFSR_71 gnd vdd FILL
XFILL_28_NOR3X1_37 gnd vdd FILL
XFILL_0_AOI21X1_11 gnd vdd FILL
XFILL_28_NOR3X1_48 gnd vdd FILL
XFILL_78_DFFSR_204 gnd vdd FILL
XFILL_18_DFFSR_82 gnd vdd FILL
XFILL_78_DFFSR_215 gnd vdd FILL
XOAI22X1_8 INVX1_86/Y OAI22X1_8/B INVX1_97/Y OAI22X1_8/D gnd OAI22X1_8/Y vdd OAI22X1
XFILL_18_DFFSR_93 gnd vdd FILL
XFILL_0_AOI21X1_22 gnd vdd FILL
XFILL_0_AOI21X1_33 gnd vdd FILL
XFILL_78_DFFSR_226 gnd vdd FILL
XFILL_0_AOI21X1_44 gnd vdd FILL
XFILL_78_DFFSR_237 gnd vdd FILL
XFILL_78_DFFSR_248 gnd vdd FILL
XFILL_29_NOR3X1_1 gnd vdd FILL
XFILL_0_AOI21X1_55 gnd vdd FILL
XFILL_13_DFFSR_170 gnd vdd FILL
XFILL_0_AOI21X1_66 gnd vdd FILL
XFILL_2_CLKBUF1_2 gnd vdd FILL
XFILL_78_DFFSR_259 gnd vdd FILL
XFILL_10_OAI22X1_13 gnd vdd FILL
XFILL_10_OAI22X1_24 gnd vdd FILL
XFILL_13_DFFSR_181 gnd vdd FILL
XFILL_10_OAI22X1_35 gnd vdd FILL
XFILL_0_AOI21X1_77 gnd vdd FILL
XFILL_13_DFFSR_192 gnd vdd FILL
XFILL_10_OAI22X1_46 gnd vdd FILL
XFILL_58_DFFSR_70 gnd vdd FILL
XFILL_58_DFFSR_81 gnd vdd FILL
XFILL_14_OAI21X1_15 gnd vdd FILL
XFILL_3_NOR2X1_110 gnd vdd FILL
XFILL_58_DFFSR_92 gnd vdd FILL
XFILL_14_OAI21X1_26 gnd vdd FILL
XFILL_3_NOR2X1_121 gnd vdd FILL
XFILL_3_NOR2X1_132 gnd vdd FILL
XFILL_3_NOR2X1_143 gnd vdd FILL
XFILL_14_OAI21X1_37 gnd vdd FILL
XFILL_59_5_0 gnd vdd FILL
XFILL_14_OAI21X1_48 gnd vdd FILL
XFILL_3_NOR2X1_154 gnd vdd FILL
XFILL_6_CLKBUF1_1 gnd vdd FILL
XFILL_3_NOR2X1_2 gnd vdd FILL
XFILL_17_DFFSR_180 gnd vdd FILL
XFILL_3_NOR2X1_165 gnd vdd FILL
XFILL_6_2_2 gnd vdd FILL
XFILL_3_NOR2X1_176 gnd vdd FILL
XFILL_17_DFFSR_191 gnd vdd FILL
XFILL_3_NOR2X1_187 gnd vdd FILL
XFILL_3_NOR2X1_198 gnd vdd FILL
XFILL_27_DFFSR_80 gnd vdd FILL
XFILL_27_DFFSR_91 gnd vdd FILL
XFILL_20_MUX2X1_101 gnd vdd FILL
XFILL_20_MUX2X1_112 gnd vdd FILL
XFILL_20_MUX2X1_123 gnd vdd FILL
XFILL_20_MUX2X1_134 gnd vdd FILL
XFILL_20_MUX2X1_145 gnd vdd FILL
XFILL_42_4_0 gnd vdd FILL
XFILL_67_DFFSR_90 gnd vdd FILL
XFILL_14_1_2 gnd vdd FILL
XFILL_20_MUX2X1_156 gnd vdd FILL
XFILL_63_DFFSR_270 gnd vdd FILL
XFILL_20_MUX2X1_167 gnd vdd FILL
XFILL_3_MUX2X1_105 gnd vdd FILL
XFILL_3_MUX2X1_116 gnd vdd FILL
XFILL_20_MUX2X1_178 gnd vdd FILL
XFILL_20_MUX2X1_189 gnd vdd FILL
XFILL_3_MUX2X1_127 gnd vdd FILL
XFILL_3_MUX2X1_138 gnd vdd FILL
XFILL_3_MUX2X1_149 gnd vdd FILL
XFILL_0_OAI22X1_30 gnd vdd FILL
XFILL_0_OAI22X1_41 gnd vdd FILL
XFILL_19_INVX8_4 gnd vdd FILL
XFILL_4_OAI21X1_10 gnd vdd FILL
XFILL_4_OAI21X1_21 gnd vdd FILL
XFILL_41_DFFSR_205 gnd vdd FILL
XFILL_4_OAI21X1_32 gnd vdd FILL
XFILL_0_NOR2X1_20 gnd vdd FILL
XFILL_4_OAI21X1_43 gnd vdd FILL
XFILL_3_OAI21X1_6 gnd vdd FILL
XFILL_0_NOR2X1_31 gnd vdd FILL
XFILL_41_DFFSR_216 gnd vdd FILL
XFILL_0_NOR2X1_42 gnd vdd FILL
XFILL_41_DFFSR_227 gnd vdd FILL
XFILL_0_NOR2X1_53 gnd vdd FILL
XFILL_41_DFFSR_238 gnd vdd FILL
XFILL_41_DFFSR_249 gnd vdd FILL
XFILL_0_NOR2X1_64 gnd vdd FILL
XFILL_0_NOR2X1_75 gnd vdd FILL
XFILL_0_NOR2X1_86 gnd vdd FILL
XFILL_0_NOR2X1_97 gnd vdd FILL
XFILL_45_DFFSR_204 gnd vdd FILL
XFILL_45_DFFSR_215 gnd vdd FILL
XFILL_23_DFFSR_6 gnd vdd FILL
XFILL_7_OAI21X1_5 gnd vdd FILL
XFILL_4_NOR2X1_30 gnd vdd FILL
XFILL_4_NOR2X1_41 gnd vdd FILL
XFILL_45_DFFSR_226 gnd vdd FILL
XFILL_80_DFFSR_7 gnd vdd FILL
XFILL_4_NOR2X1_52 gnd vdd FILL
XFILL_45_DFFSR_237 gnd vdd FILL
XFILL_45_DFFSR_248 gnd vdd FILL
XFILL_4_NOR2X1_63 gnd vdd FILL
XFILL_45_DFFSR_259 gnd vdd FILL
XFILL_4_NOR2X1_74 gnd vdd FILL
XFILL_4_NOR2X1_85 gnd vdd FILL
XFILL_4_NOR2X1_96 gnd vdd FILL
XFILL_72_DFFSR_104 gnd vdd FILL
XFILL_49_DFFSR_203 gnd vdd FILL
XFILL_72_DFFSR_115 gnd vdd FILL
XFILL_49_DFFSR_214 gnd vdd FILL
XFILL_72_DFFSR_126 gnd vdd FILL
XFILL_49_DFFSR_225 gnd vdd FILL
XFILL_72_DFFSR_137 gnd vdd FILL
XFILL_8_NOR2X1_40 gnd vdd FILL
XFILL_12_OAI22X1_2 gnd vdd FILL
XFILL_72_DFFSR_148 gnd vdd FILL
XFILL_8_NOR2X1_51 gnd vdd FILL
XFILL_49_DFFSR_236 gnd vdd FILL
XFILL_8_NOR2X1_62 gnd vdd FILL
XFILL_49_DFFSR_247 gnd vdd FILL
XFILL_49_DFFSR_258 gnd vdd FILL
XFILL_72_DFFSR_159 gnd vdd FILL
XFILL_49_DFFSR_269 gnd vdd FILL
XFILL_8_NOR2X1_73 gnd vdd FILL
XFILL_8_NOR2X1_84 gnd vdd FILL
XFILL_8_NOR2X1_95 gnd vdd FILL
XFILL_76_DFFSR_103 gnd vdd FILL
XFILL_64_0_2 gnd vdd FILL
XFILL_76_DFFSR_114 gnd vdd FILL
XFILL_6_NAND3X1_19 gnd vdd FILL
XFILL_76_DFFSR_125 gnd vdd FILL
XFILL_76_DFFSR_136 gnd vdd FILL
XFILL_16_OAI22X1_1 gnd vdd FILL
XFILL_76_DFFSR_147 gnd vdd FILL
XFILL_76_DFFSR_158 gnd vdd FILL
XFILL_76_DFFSR_169 gnd vdd FILL
XFILL_6_BUFX4_19 gnd vdd FILL
XFILL_33_4_0 gnd vdd FILL
XFILL_26_2 gnd vdd FILL
XFILL_19_1 gnd vdd FILL
XFILL_30_DFFSR_270 gnd vdd FILL
XFILL_0_NAND2X1_8 gnd vdd FILL
XFILL_4_NAND2X1_7 gnd vdd FILL
XFILL_0_MUX2X1_60 gnd vdd FILL
XFILL_0_MUX2X1_71 gnd vdd FILL
XFILL_0_MUX2X1_82 gnd vdd FILL
XFILL_0_MUX2X1_93 gnd vdd FILL
XFILL_13_AND2X2_7 gnd vdd FILL
XFILL_61_DFFSR_180 gnd vdd FILL
XFILL_61_DFFSR_191 gnd vdd FILL
XFILL_8_NAND2X1_6 gnd vdd FILL
XFILL_12_DFFSR_204 gnd vdd FILL
XFILL_12_DFFSR_215 gnd vdd FILL
XFILL_12_DFFSR_226 gnd vdd FILL
XFILL_12_DFFSR_237 gnd vdd FILL
XFILL_4_MUX2X1_70 gnd vdd FILL
XFILL_4_MUX2X1_81 gnd vdd FILL
XFILL_12_DFFSR_248 gnd vdd FILL
XFILL_4_MUX2X1_92 gnd vdd FILL
XFILL_12_DFFSR_259 gnd vdd FILL
XFILL_65_DFFSR_190 gnd vdd FILL
XFILL_10_BUFX4_13 gnd vdd FILL
XFILL_16_DFFSR_203 gnd vdd FILL
XFILL_13_NAND3X1_3 gnd vdd FILL
XFILL_10_BUFX4_24 gnd vdd FILL
XFILL_16_DFFSR_214 gnd vdd FILL
XFILL_10_BUFX4_35 gnd vdd FILL
XFILL_10_BUFX4_46 gnd vdd FILL
XFILL_16_DFFSR_225 gnd vdd FILL
XFILL_16_DFFSR_236 gnd vdd FILL
XFILL_8_MUX2X1_80 gnd vdd FILL
XFILL_10_BUFX4_57 gnd vdd FILL
XFILL_16_DFFSR_247 gnd vdd FILL
XFILL_10_BUFX4_68 gnd vdd FILL
XFILL_7_BUFX4_9 gnd vdd FILL
XFILL_8_MUX2X1_91 gnd vdd FILL
XFILL_16_DFFSR_258 gnd vdd FILL
XFILL_55_0_2 gnd vdd FILL
XFILL_16_DFFSR_269 gnd vdd FILL
XFILL_10_BUFX4_79 gnd vdd FILL
XFILL_43_DFFSR_103 gnd vdd FILL
XFILL_43_DFFSR_114 gnd vdd FILL
XFILL_43_DFFSR_125 gnd vdd FILL
XFILL_43_DFFSR_136 gnd vdd FILL
XFILL_43_DFFSR_147 gnd vdd FILL
XFILL_43_DFFSR_158 gnd vdd FILL
XFILL_24_4_0 gnd vdd FILL
XFILL_43_DFFSR_169 gnd vdd FILL
XFILL_47_DFFSR_102 gnd vdd FILL
XFILL_47_DFFSR_113 gnd vdd FILL
XFILL_47_DFFSR_124 gnd vdd FILL
XFILL_6_NOR2X1_109 gnd vdd FILL
XFILL_47_DFFSR_135 gnd vdd FILL
XFILL_47_DFFSR_146 gnd vdd FILL
XFILL_12_NAND3X1_11 gnd vdd FILL
XFILL_47_DFFSR_157 gnd vdd FILL
XFILL_12_NAND3X1_22 gnd vdd FILL
XFILL_47_DFFSR_168 gnd vdd FILL
XFILL_12_NAND3X1_33 gnd vdd FILL
XFILL_47_DFFSR_179 gnd vdd FILL
XFILL_20_MUX2X1_90 gnd vdd FILL
XFILL_12_NAND3X1_44 gnd vdd FILL
XFILL_4_INVX1_14 gnd vdd FILL
XFILL_12_NAND3X1_55 gnd vdd FILL
XFILL_4_INVX1_25 gnd vdd FILL
XFILL_32_CLKBUF1_11 gnd vdd FILL
XFILL_12_NAND3X1_66 gnd vdd FILL
XFILL_4_INVX1_36 gnd vdd FILL
XFILL_12_NAND3X1_77 gnd vdd FILL
XFILL_32_CLKBUF1_22 gnd vdd FILL
XFILL_4_INVX1_47 gnd vdd FILL
XFILL_5_AND2X2_6 gnd vdd FILL
XFILL_12_NAND3X1_88 gnd vdd FILL
XFILL_32_CLKBUF1_33 gnd vdd FILL
XFILL_4_INVX1_58 gnd vdd FILL
XFILL_12_NAND3X1_99 gnd vdd FILL
XFILL_4_INVX1_69 gnd vdd FILL
XFILL_3_BUFX2_5 gnd vdd FILL
XFILL_13_AOI22X1_8 gnd vdd FILL
XFILL_17_AOI22X1_7 gnd vdd FILL
XFILL_2_BUFX4_12 gnd vdd FILL
XFILL_62_DFFSR_4 gnd vdd FILL
XFILL_2_BUFX4_23 gnd vdd FILL
XFILL_2_BUFX4_34 gnd vdd FILL
XFILL_2_BUFX4_45 gnd vdd FILL
XFILL_19_DFFSR_16 gnd vdd FILL
XFILL_2_BUFX4_56 gnd vdd FILL
XFILL_1_OR2X2_1 gnd vdd FILL
XFILL_7_5_0 gnd vdd FILL
XFILL_19_DFFSR_27 gnd vdd FILL
XFILL_2_BUFX4_67 gnd vdd FILL
XFILL_19_DFFSR_38 gnd vdd FILL
XFILL_2_BUFX4_78 gnd vdd FILL
XFILL_19_DFFSR_49 gnd vdd FILL
XFILL_3_OAI22X1_18 gnd vdd FILL
XFILL_2_BUFX4_89 gnd vdd FILL
XFILL_3_OAI22X1_29 gnd vdd FILL
XFILL_32_DFFSR_190 gnd vdd FILL
XFILL_59_DFFSR_15 gnd vdd FILL
XFILL_16_AOI22X1_11 gnd vdd FILL
XFILL_59_DFFSR_26 gnd vdd FILL
XFILL_46_0_2 gnd vdd FILL
XFILL_59_DFFSR_37 gnd vdd FILL
XFILL_59_DFFSR_48 gnd vdd FILL
XFILL_59_DFFSR_59 gnd vdd FILL
XFILL_2_NAND3X1_50 gnd vdd FILL
XFILL_2_NAND3X1_61 gnd vdd FILL
XFILL_2_NAND3X1_72 gnd vdd FILL
XFILL_2_NAND3X1_83 gnd vdd FILL
XFILL_6_NAND2X1_30 gnd vdd FILL
XFILL_2_NAND3X1_94 gnd vdd FILL
XFILL_10_DFFSR_103 gnd vdd FILL
XFILL_6_NAND2X1_41 gnd vdd FILL
XFILL_6_NAND2X1_52 gnd vdd FILL
XFILL_10_DFFSR_114 gnd vdd FILL
XFILL_15_4_0 gnd vdd FILL
XFILL_27_DFFSR_7 gnd vdd FILL
XFILL_6_NAND2X1_63 gnd vdd FILL
XFILL_10_DFFSR_125 gnd vdd FILL
XFILL_10_DFFSR_136 gnd vdd FILL
XFILL_6_NAND2X1_74 gnd vdd FILL
XFILL_84_DFFSR_8 gnd vdd FILL
XFILL_28_DFFSR_14 gnd vdd FILL
XMUX2X1_1 MUX2X1_1/A MUX2X1_1/B MUX2X1_1/S gnd MUX2X1_1/Y vdd MUX2X1
XFILL_28_DFFSR_25 gnd vdd FILL
XFILL_6_NAND2X1_85 gnd vdd FILL
XFILL_10_DFFSR_147 gnd vdd FILL
XFILL_10_DFFSR_158 gnd vdd FILL
XFILL_6_NAND2X1_96 gnd vdd FILL
XFILL_28_DFFSR_36 gnd vdd FILL
XFILL_10_DFFSR_169 gnd vdd FILL
XFILL_3_INVX2_5 gnd vdd FILL
XFILL_28_DFFSR_47 gnd vdd FILL
XFILL_14_DFFSR_102 gnd vdd FILL
XFILL_28_DFFSR_58 gnd vdd FILL
XFILL_28_DFFSR_69 gnd vdd FILL
XFILL_14_CLKBUF1_16 gnd vdd FILL
XFILL_14_DFFSR_113 gnd vdd FILL
XFILL_14_DFFSR_124 gnd vdd FILL
XFILL_14_CLKBUF1_27 gnd vdd FILL
XFILL_14_CLKBUF1_38 gnd vdd FILL
XFILL_14_DFFSR_135 gnd vdd FILL
XFILL_14_DFFSR_146 gnd vdd FILL
XFILL_68_DFFSR_13 gnd vdd FILL
XFILL_68_DFFSR_24 gnd vdd FILL
XFILL_14_DFFSR_157 gnd vdd FILL
XFILL_68_DFFSR_35 gnd vdd FILL
XFILL_14_DFFSR_168 gnd vdd FILL
XFILL_14_DFFSR_179 gnd vdd FILL
XFILL_68_DFFSR_46 gnd vdd FILL
XFILL_18_DFFSR_101 gnd vdd FILL
XFILL_68_DFFSR_57 gnd vdd FILL
XFILL_68_DFFSR_68 gnd vdd FILL
XFILL_68_DFFSR_79 gnd vdd FILL
XFILL_18_DFFSR_112 gnd vdd FILL
XFILL_1_INVX1_3 gnd vdd FILL
XFILL_18_DFFSR_123 gnd vdd FILL
XFILL_18_DFFSR_134 gnd vdd FILL
XFILL_18_DFFSR_145 gnd vdd FILL
XFILL_18_DFFSR_156 gnd vdd FILL
XCLKBUF1_2 BUFX4_73/Y gnd DFFSR_2/CLK vdd CLKBUF1
XFILL_18_DFFSR_167 gnd vdd FILL
XFILL_18_DFFSR_178 gnd vdd FILL
XFILL_10_NOR3X1_14 gnd vdd FILL
XFILL_37_DFFSR_12 gnd vdd FILL
XFILL_18_DFFSR_189 gnd vdd FILL
XFILL_10_NOR3X1_25 gnd vdd FILL
XFILL_37_DFFSR_23 gnd vdd FILL
XFILL_10_NOR3X1_36 gnd vdd FILL
XFILL_37_DFFSR_34 gnd vdd FILL
XFILL_10_NOR3X1_47 gnd vdd FILL
XFILL_60_DFFSR_203 gnd vdd FILL
XFILL_37_DFFSR_45 gnd vdd FILL
XFILL_60_DFFSR_214 gnd vdd FILL
XFILL_37_DFFSR_56 gnd vdd FILL
XFILL_37_DFFSR_67 gnd vdd FILL
XFILL_3_BUFX4_105 gnd vdd FILL
XFILL_60_DFFSR_225 gnd vdd FILL
XFILL_37_DFFSR_78 gnd vdd FILL
XFILL_60_DFFSR_236 gnd vdd FILL
XFILL_37_DFFSR_89 gnd vdd FILL
XFILL_60_DFFSR_247 gnd vdd FILL
XFILL_14_NOR3X1_13 gnd vdd FILL
XFILL_60_DFFSR_258 gnd vdd FILL
XFILL_77_DFFSR_11 gnd vdd FILL
XFILL_14_NOR3X1_24 gnd vdd FILL
XFILL_60_DFFSR_269 gnd vdd FILL
XFILL_77_DFFSR_22 gnd vdd FILL
XFILL_14_NOR3X1_35 gnd vdd FILL
XFILL_77_DFFSR_33 gnd vdd FILL
XFILL_64_DFFSR_202 gnd vdd FILL
XFILL_14_NOR3X1_46 gnd vdd FILL
XFILL_77_DFFSR_44 gnd vdd FILL
XFILL_77_DFFSR_55 gnd vdd FILL
XFILL_64_DFFSR_213 gnd vdd FILL
XFILL_21_CLKBUF1_40 gnd vdd FILL
XFILL_64_DFFSR_224 gnd vdd FILL
XFILL_7_BUFX4_104 gnd vdd FILL
XFILL_77_DFFSR_66 gnd vdd FILL
XFILL_77_DFFSR_77 gnd vdd FILL
XFILL_64_DFFSR_235 gnd vdd FILL
XFILL_65_3_0 gnd vdd FILL
XFILL_77_DFFSR_88 gnd vdd FILL
XFILL_64_DFFSR_246 gnd vdd FILL
XFILL_4_CLKBUF1_11 gnd vdd FILL
XFILL_77_DFFSR_99 gnd vdd FILL
XFILL_37_0_2 gnd vdd FILL
XFILL_18_NOR3X1_12 gnd vdd FILL
XFILL_64_DFFSR_257 gnd vdd FILL
XFILL_4_CLKBUF1_22 gnd vdd FILL
XFILL_64_DFFSR_268 gnd vdd FILL
XFILL_18_NOR3X1_23 gnd vdd FILL
XFILL_0_INVX1_40 gnd vdd FILL
XFILL_18_NOR3X1_34 gnd vdd FILL
XNOR2X1_200 DFFSR_7/Q NOR2X1_202/B gnd NOR2X1_200/Y vdd NOR2X1
XFILL_4_CLKBUF1_33 gnd vdd FILL
XFILL_0_INVX1_51 gnd vdd FILL
XFILL_68_DFFSR_201 gnd vdd FILL
XFILL_0_INVX1_62 gnd vdd FILL
XFILL_18_NOR3X1_45 gnd vdd FILL
XFILL_68_DFFSR_212 gnd vdd FILL
XFILL_46_DFFSR_10 gnd vdd FILL
XFILL_0_INVX1_73 gnd vdd FILL
XFILL_12_MUX2X1_107 gnd vdd FILL
XFILL_0_INVX1_84 gnd vdd FILL
XFILL_12_MUX2X1_118 gnd vdd FILL
XFILL_68_DFFSR_223 gnd vdd FILL
XFILL_12_MUX2X1_129 gnd vdd FILL
XFILL_46_DFFSR_21 gnd vdd FILL
XFILL_0_INVX1_95 gnd vdd FILL
XFILL_68_DFFSR_234 gnd vdd FILL
XFILL_46_DFFSR_32 gnd vdd FILL
XFILL_46_DFFSR_43 gnd vdd FILL
XFILL_68_DFFSR_245 gnd vdd FILL
XFILL_17_NOR3X1_7 gnd vdd FILL
XFILL_68_DFFSR_256 gnd vdd FILL
XFILL_46_DFFSR_54 gnd vdd FILL
XFILL_68_DFFSR_267 gnd vdd FILL
XFILL_46_DFFSR_65 gnd vdd FILL
XFILL_23_CLKBUF1_8 gnd vdd FILL
XFILL_46_DFFSR_76 gnd vdd FILL
XFILL_46_DFFSR_87 gnd vdd FILL
XFILL_1_NOR2X1_18 gnd vdd FILL
XFILL_46_DFFSR_98 gnd vdd FILL
XFILL_13_OAI21X1_12 gnd vdd FILL
XFILL_1_NOR2X1_29 gnd vdd FILL
XFILL_86_DFFSR_20 gnd vdd FILL
XFILL_13_OAI21X1_23 gnd vdd FILL
XFILL_13_OAI21X1_34 gnd vdd FILL
XFILL_2_NOR2X1_140 gnd vdd FILL
XFILL_86_DFFSR_31 gnd vdd FILL
XFILL_2_NOR2X1_151 gnd vdd FILL
XFILL_86_DFFSR_42 gnd vdd FILL
XFILL_13_OAI21X1_45 gnd vdd FILL
XFILL_2_NOR2X1_162 gnd vdd FILL
XFILL_86_DFFSR_53 gnd vdd FILL
XFILL_15_DFFSR_20 gnd vdd FILL
XFILL_86_DFFSR_64 gnd vdd FILL
XFILL_27_CLKBUF1_7 gnd vdd FILL
XFILL_2_NOR2X1_173 gnd vdd FILL
XFILL_86_DFFSR_75 gnd vdd FILL
XFILL_2_NOR2X1_184 gnd vdd FILL
XFILL_15_DFFSR_31 gnd vdd FILL
XFILL_86_DFFSR_86 gnd vdd FILL
XFILL_15_DFFSR_42 gnd vdd FILL
XFILL_2_NOR2X1_195 gnd vdd FILL
XFILL_15_DFFSR_53 gnd vdd FILL
XFILL_86_DFFSR_97 gnd vdd FILL
XFILL_5_NOR2X1_17 gnd vdd FILL
XFILL_5_NOR2X1_28 gnd vdd FILL
XFILL_15_DFFSR_64 gnd vdd FILL
XFILL_15_DFFSR_75 gnd vdd FILL
XFILL_5_NOR2X1_39 gnd vdd FILL
XFILL_15_DFFSR_86 gnd vdd FILL
XFILL_15_DFFSR_97 gnd vdd FILL
XFILL_55_DFFSR_30 gnd vdd FILL
XFILL_26_NOR3X1_5 gnd vdd FILL
XFILL_55_DFFSR_41 gnd vdd FILL
XFILL_9_NOR2X1_16 gnd vdd FILL
XFILL_55_DFFSR_52 gnd vdd FILL
XFILL_55_DFFSR_63 gnd vdd FILL
XFILL_9_NOR2X1_27 gnd vdd FILL
XFILL_55_DFFSR_74 gnd vdd FILL
XFILL_9_NOR2X1_38 gnd vdd FILL
XFILL_55_DFFSR_85 gnd vdd FILL
XFILL_9_NOR2X1_49 gnd vdd FILL
XFILL_55_DFFSR_96 gnd vdd FILL
XFILL_2_MUX2X1_102 gnd vdd FILL
XFILL_2_MUX2X1_113 gnd vdd FILL
XFILL_0_NOR2X1_6 gnd vdd FILL
XFILL_2_MUX2X1_124 gnd vdd FILL
XFILL_44_DFFSR_1 gnd vdd FILL
XFILL_2_MUX2X1_135 gnd vdd FILL
XFILL_2_MUX2X1_146 gnd vdd FILL
XFILL_24_DFFSR_40 gnd vdd FILL
XFILL_2_MUX2X1_157 gnd vdd FILL
XFILL_2_MUX2X1_168 gnd vdd FILL
XFILL_24_DFFSR_51 gnd vdd FILL
XFILL_2_MUX2X1_179 gnd vdd FILL
XFILL_24_DFFSR_62 gnd vdd FILL
XFILL_24_DFFSR_73 gnd vdd FILL
XFILL_24_DFFSR_84 gnd vdd FILL
XFILL_24_DFFSR_95 gnd vdd FILL
XFILL_31_DFFSR_202 gnd vdd FILL
XFILL_56_3_0 gnd vdd FILL
XFILL_9_NOR3X1_6 gnd vdd FILL
XFILL_31_DFFSR_213 gnd vdd FILL
XFILL_3_OAI21X1_40 gnd vdd FILL
XFILL_3_0_2 gnd vdd FILL
XFILL_28_0_2 gnd vdd FILL
XFILL_7_BUFX2_6 gnd vdd FILL
XFILL_31_DFFSR_224 gnd vdd FILL
XFILL_31_DFFSR_235 gnd vdd FILL
XFILL_64_DFFSR_50 gnd vdd FILL
XFILL_31_DFFSR_246 gnd vdd FILL
XFILL_0_DFFSR_270 gnd vdd FILL
XFILL_31_DFFSR_257 gnd vdd FILL
XFILL_64_DFFSR_61 gnd vdd FILL
XFILL_31_DFFSR_268 gnd vdd FILL
XFILL_64_DFFSR_72 gnd vdd FILL
XFILL_64_DFFSR_83 gnd vdd FILL
XFILL_64_DFFSR_94 gnd vdd FILL
XFILL_35_DFFSR_201 gnd vdd FILL
XFILL_35_DFFSR_212 gnd vdd FILL
XFILL_35_DFFSR_223 gnd vdd FILL
XFILL_35_DFFSR_234 gnd vdd FILL
XFILL_7_DFFSR_30 gnd vdd FILL
XFILL_35_DFFSR_245 gnd vdd FILL
XFILL_7_DFFSR_41 gnd vdd FILL
XFILL_66_DFFSR_5 gnd vdd FILL
XFILL_35_DFFSR_256 gnd vdd FILL
XFILL_35_DFFSR_267 gnd vdd FILL
XFILL_7_DFFSR_52 gnd vdd FILL
XFILL_7_DFFSR_63 gnd vdd FILL
XFILL_40_7_1 gnd vdd FILL
XFILL_1_MUX2X1_14 gnd vdd FILL
XFILL_1_MUX2X1_25 gnd vdd FILL
XFILL_62_DFFSR_101 gnd vdd FILL
XFILL_7_DFFSR_74 gnd vdd FILL
XFILL_39_DFFSR_200 gnd vdd FILL
XFILL_7_DFFSR_85 gnd vdd FILL
XFILL_33_DFFSR_60 gnd vdd FILL
XFILL_1_MUX2X1_36 gnd vdd FILL
XINVX8_4 din[0] gnd INVX8_4/Y vdd INVX8
XFILL_39_DFFSR_211 gnd vdd FILL
XFILL_1_MUX2X1_47 gnd vdd FILL
XFILL_7_DFFSR_96 gnd vdd FILL
XFILL_62_DFFSR_112 gnd vdd FILL
XFILL_39_DFFSR_222 gnd vdd FILL
XFILL_1_MUX2X1_58 gnd vdd FILL
XFILL_33_DFFSR_71 gnd vdd FILL
XFILL_62_DFFSR_123 gnd vdd FILL
XFILL_33_DFFSR_82 gnd vdd FILL
XFILL_62_DFFSR_134 gnd vdd FILL
XFILL_39_DFFSR_233 gnd vdd FILL
XFILL_1_MUX2X1_69 gnd vdd FILL
XFILL_33_DFFSR_93 gnd vdd FILL
XFILL_62_DFFSR_145 gnd vdd FILL
XFILL_62_DFFSR_156 gnd vdd FILL
XFILL_39_DFFSR_244 gnd vdd FILL
XFILL_39_DFFSR_255 gnd vdd FILL
XFILL_5_MUX2X1_13 gnd vdd FILL
XFILL_62_DFFSR_167 gnd vdd FILL
XFILL_39_DFFSR_266 gnd vdd FILL
XFILL_62_DFFSR_178 gnd vdd FILL
XFILL_66_DFFSR_100 gnd vdd FILL
XFILL_62_DFFSR_189 gnd vdd FILL
XFILL_5_MUX2X1_24 gnd vdd FILL
XFILL_5_MUX2X1_35 gnd vdd FILL
XFILL_66_DFFSR_111 gnd vdd FILL
XFILL_73_DFFSR_70 gnd vdd FILL
XFILL_5_MUX2X1_46 gnd vdd FILL
XFILL_5_NAND3X1_16 gnd vdd FILL
XFILL_5_MUX2X1_57 gnd vdd FILL
XFILL_66_DFFSR_122 gnd vdd FILL
XFILL_66_DFFSR_133 gnd vdd FILL
XFILL_5_NAND3X1_27 gnd vdd FILL
XFILL_73_DFFSR_81 gnd vdd FILL
XFILL_73_DFFSR_92 gnd vdd FILL
XFILL_66_DFFSR_144 gnd vdd FILL
XFILL_5_MUX2X1_68 gnd vdd FILL
XFILL_5_NAND3X1_38 gnd vdd FILL
XFILL_5_MUX2X1_79 gnd vdd FILL
XFILL_66_DFFSR_155 gnd vdd FILL
XFILL_5_NAND3X1_49 gnd vdd FILL
XFILL_9_NAND2X1_18 gnd vdd FILL
XFILL_66_DFFSR_166 gnd vdd FILL
XFILL_9_MUX2X1_12 gnd vdd FILL
XFILL_66_DFFSR_177 gnd vdd FILL
XFILL_9_MUX2X1_23 gnd vdd FILL
XFILL_66_DFFSR_188 gnd vdd FILL
XFILL_9_NAND2X1_29 gnd vdd FILL
XFILL_9_MUX2X1_34 gnd vdd FILL
XFILL_66_DFFSR_199 gnd vdd FILL
XFILL_9_MUX2X1_45 gnd vdd FILL
XFILL_9_MUX2X1_56 gnd vdd FILL
XFILL_9_MUX2X1_67 gnd vdd FILL
XFILL_9_MUX2X1_78 gnd vdd FILL
XFILL_9_MUX2X1_89 gnd vdd FILL
XFILL_42_DFFSR_80 gnd vdd FILL
XFILL_19_MUX2X1_160 gnd vdd FILL
XFILL_42_DFFSR_91 gnd vdd FILL
XBUFX4_13 BUFX4_51/Y gnd BUFX4_13/Y vdd BUFX4
XFILL_10_NOR2X1_80 gnd vdd FILL
XFILL_19_MUX2X1_171 gnd vdd FILL
XBUFX4_24 BUFX4_51/Y gnd DFFSR_49/R vdd BUFX4
XFILL_19_MUX2X1_182 gnd vdd FILL
XFILL_10_NOR2X1_91 gnd vdd FILL
XBUFX4_35 BUFX4_54/A gnd DFFSR_5/R vdd BUFX4
XFILL_19_MUX2X1_193 gnd vdd FILL
XBUFX4_46 BUFX4_51/Y gnd DFFSR_45/R vdd BUFX4
XBUFX4_57 BUFX4_60/A gnd BUFX4_57/Y vdd BUFX4
XBUFX4_68 INVX8_1/Y gnd BUFX4_68/Y vdd BUFX4
XFILL_47_3_0 gnd vdd FILL
XBUFX4_79 INVX8_4/Y gnd MUX2X1_8/A vdd BUFX4
XFILL_82_DFFSR_90 gnd vdd FILL
XFILL_19_0_2 gnd vdd FILL
XFILL_21_MUX2X1_11 gnd vdd FILL
XFILL_21_MUX2X1_22 gnd vdd FILL
XFILL_5_INVX1_4 gnd vdd FILL
XFILL_21_MUX2X1_33 gnd vdd FILL
XFILL_11_DFFSR_90 gnd vdd FILL
XFILL_21_MUX2X1_44 gnd vdd FILL
XFILL_21_MUX2X1_55 gnd vdd FILL
XFILL_21_MUX2X1_66 gnd vdd FILL
XFILL_21_MUX2X1_77 gnd vdd FILL
XFILL_21_MUX2X1_88 gnd vdd FILL
XFILL_21_MUX2X1_99 gnd vdd FILL
XFILL_31_7_1 gnd vdd FILL
XFILL_10_5 gnd vdd FILL
XFILL_30_2_0 gnd vdd FILL
XFILL_24_CLKBUF1_17 gnd vdd FILL
XFILL_24_CLKBUF1_28 gnd vdd FILL
XFILL_24_CLKBUF1_39 gnd vdd FILL
XFILL_33_DFFSR_100 gnd vdd FILL
XFILL_33_DFFSR_111 gnd vdd FILL
XFILL_10_NAND2X1_2 gnd vdd FILL
XFILL_2_AOI21X1_18 gnd vdd FILL
XFILL_33_DFFSR_122 gnd vdd FILL
XFILL_33_DFFSR_133 gnd vdd FILL
XFILL_33_DFFSR_144 gnd vdd FILL
XFILL_2_AOI21X1_29 gnd vdd FILL
XFILL_33_DFFSR_155 gnd vdd FILL
XFILL_33_DFFSR_166 gnd vdd FILL
XFILL_33_DFFSR_177 gnd vdd FILL
XFILL_2_DFFSR_190 gnd vdd FILL
XFILL_33_DFFSR_188 gnd vdd FILL
XFILL_37_DFFSR_110 gnd vdd FILL
XFILL_33_DFFSR_199 gnd vdd FILL
XFILL_5_NOR2X1_106 gnd vdd FILL
XFILL_37_DFFSR_121 gnd vdd FILL
XFILL_37_DFFSR_132 gnd vdd FILL
XFILL_5_NOR2X1_117 gnd vdd FILL
XFILL_37_DFFSR_143 gnd vdd FILL
XFILL_5_NOR2X1_128 gnd vdd FILL
XFILL_37_DFFSR_154 gnd vdd FILL
XFILL_5_NOR2X1_139 gnd vdd FILL
XFILL_37_DFFSR_165 gnd vdd FILL
XFILL_11_NAND3X1_30 gnd vdd FILL
XFILL_11_NAND3X1_41 gnd vdd FILL
XFILL_37_DFFSR_176 gnd vdd FILL
XFILL_37_DFFSR_187 gnd vdd FILL
XFILL_11_NAND3X1_52 gnd vdd FILL
XFILL_37_DFFSR_198 gnd vdd FILL
XFILL_11_NAND3X1_63 gnd vdd FILL
XFILL_11_NAND3X1_74 gnd vdd FILL
XFILL_11_NAND3X1_85 gnd vdd FILL
XFILL_38_3_0 gnd vdd FILL
XFILL_31_CLKBUF1_30 gnd vdd FILL
XFILL_31_CLKBUF1_41 gnd vdd FILL
XFILL_11_NAND3X1_96 gnd vdd FILL
XFILL_83_DFFSR_200 gnd vdd FILL
XFILL_22_MUX2X1_108 gnd vdd FILL
XFILL_83_DFFSR_211 gnd vdd FILL
XFILL_22_MUX2X1_119 gnd vdd FILL
XFILL_83_DFFSR_222 gnd vdd FILL
XFILL_10_DFFSR_4 gnd vdd FILL
XFILL_10_AOI21X1_7 gnd vdd FILL
XFILL_83_DFFSR_233 gnd vdd FILL
XFILL_83_DFFSR_244 gnd vdd FILL
XFILL_83_DFFSR_255 gnd vdd FILL
XFILL_83_DFFSR_266 gnd vdd FILL
XFILL_22_7_1 gnd vdd FILL
XFILL_48_DFFSR_2 gnd vdd FILL
XFILL_1_INVX1_18 gnd vdd FILL
XFILL_21_2_0 gnd vdd FILL
XFILL_87_DFFSR_210 gnd vdd FILL
XFILL_1_INVX1_29 gnd vdd FILL
XFILL_87_DFFSR_221 gnd vdd FILL
XFILL_14_AOI21X1_6 gnd vdd FILL
XFILL_2_OAI22X1_15 gnd vdd FILL
XFILL_87_DFFSR_232 gnd vdd FILL
XFILL_2_OAI22X1_26 gnd vdd FILL
XFILL_87_DFFSR_243 gnd vdd FILL
XFILL_87_DFFSR_254 gnd vdd FILL
XFILL_2_OAI22X1_37 gnd vdd FILL
XFILL_87_DFFSR_265 gnd vdd FILL
XFILL_2_OAI22X1_48 gnd vdd FILL
XFILL_6_OAI21X1_17 gnd vdd FILL
XFILL_6_OAI21X1_28 gnd vdd FILL
XFILL_6_OAI21X1_39 gnd vdd FILL
XFILL_3_INVX1_160 gnd vdd FILL
XFILL_3_INVX1_171 gnd vdd FILL
XFILL_3_INVX1_182 gnd vdd FILL
XFILL_3_INVX1_193 gnd vdd FILL
XFILL_1_NAND3X1_80 gnd vdd FILL
XFILL_1_NAND3X1_91 gnd vdd FILL
XFILL_32_DFFSR_8 gnd vdd FILL
XFILL_5_NAND2X1_60 gnd vdd FILL
XFILL_5_NAND2X1_71 gnd vdd FILL
XFILL_5_NAND2X1_82 gnd vdd FILL
XFILL_7_INVX1_170 gnd vdd FILL
XFILL_5_NAND2X1_93 gnd vdd FILL
XFILL_7_INVX1_181 gnd vdd FILL
XFILL_7_INVX1_192 gnd vdd FILL
XFILL_13_CLKBUF1_13 gnd vdd FILL
XFILL_13_CLKBUF1_24 gnd vdd FILL
XFILL_56_DFFSR_19 gnd vdd FILL
XFILL_13_CLKBUF1_35 gnd vdd FILL
XFILL_29_3_0 gnd vdd FILL
XFILL_4_3_0 gnd vdd FILL
XFILL_11_NOR2X1_120 gnd vdd FILL
XFILL_11_NOR2X1_131 gnd vdd FILL
XFILL_25_DFFSR_18 gnd vdd FILL
XFILL_11_NOR2X1_142 gnd vdd FILL
XFILL_25_DFFSR_29 gnd vdd FILL
XFILL_11_NOR2X1_153 gnd vdd FILL
XFILL_11_NOR2X1_164 gnd vdd FILL
XFILL_50_DFFSR_200 gnd vdd FILL
XFILL_11_NOR2X1_175 gnd vdd FILL
XFILL_50_DFFSR_211 gnd vdd FILL
XFILL_11_NOR2X1_186 gnd vdd FILL
XFILL_50_DFFSR_222 gnd vdd FILL
XFILL_11_NOR2X1_197 gnd vdd FILL
XFILL_13_7_1 gnd vdd FILL
XFILL_50_DFFSR_233 gnd vdd FILL
XFILL_50_DFFSR_244 gnd vdd FILL
XFILL_50_DFFSR_255 gnd vdd FILL
XFILL_65_DFFSR_17 gnd vdd FILL
XFILL_12_2_0 gnd vdd FILL
XFILL_65_DFFSR_28 gnd vdd FILL
XFILL_9_AOI21X1_60 gnd vdd FILL
XFILL_50_DFFSR_266 gnd vdd FILL
XFILL_9_AOI21X1_71 gnd vdd FILL
XFILL_65_DFFSR_39 gnd vdd FILL
XFILL_19_OAI22X1_40 gnd vdd FILL
XFILL_19_OAI22X1_51 gnd vdd FILL
XFILL_54_DFFSR_210 gnd vdd FILL
XFILL_54_DFFSR_221 gnd vdd FILL
XFILL_54_DFFSR_232 gnd vdd FILL
XFILL_54_DFFSR_243 gnd vdd FILL
XFILL_54_DFFSR_254 gnd vdd FILL
XFILL_54_DFFSR_265 gnd vdd FILL
XFILL_3_CLKBUF1_30 gnd vdd FILL
XFILL_8_DFFSR_19 gnd vdd FILL
XFILL_3_CLKBUF1_41 gnd vdd FILL
XFILL_11_MUX2X1_104 gnd vdd FILL
XFILL_34_DFFSR_16 gnd vdd FILL
XFILL_81_DFFSR_110 gnd vdd FILL
XFILL_11_MUX2X1_115 gnd vdd FILL
XFILL_58_DFFSR_220 gnd vdd FILL
XFILL_34_DFFSR_27 gnd vdd FILL
XFILL_81_DFFSR_121 gnd vdd FILL
XFILL_81_DFFSR_132 gnd vdd FILL
XFILL_34_DFFSR_38 gnd vdd FILL
XFILL_11_MUX2X1_126 gnd vdd FILL
XFILL_58_DFFSR_231 gnd vdd FILL
XFILL_81_DFFSR_143 gnd vdd FILL
XFILL_11_MUX2X1_137 gnd vdd FILL
XFILL_34_DFFSR_49 gnd vdd FILL
XFILL_81_DFFSR_154 gnd vdd FILL
XFILL_58_DFFSR_242 gnd vdd FILL
XFILL_11_MUX2X1_148 gnd vdd FILL
XFILL_11_MUX2X1_159 gnd vdd FILL
XFILL_58_DFFSR_253 gnd vdd FILL
XFILL_81_DFFSR_165 gnd vdd FILL
XFILL_58_DFFSR_264 gnd vdd FILL
XFILL_58_DFFSR_275 gnd vdd FILL
XFILL_81_DFFSR_176 gnd vdd FILL
XFILL_13_CLKBUF1_5 gnd vdd FILL
XFILL_1_DFFSR_202 gnd vdd FILL
XFILL_81_DFFSR_187 gnd vdd FILL
XFILL_1_DFFSR_213 gnd vdd FILL
XFILL_81_DFFSR_198 gnd vdd FILL
XFILL_74_DFFSR_15 gnd vdd FILL
XFILL_1_DFFSR_224 gnd vdd FILL
XFILL_12_OAI21X1_20 gnd vdd FILL
XFILL_85_DFFSR_120 gnd vdd FILL
XFILL_74_DFFSR_26 gnd vdd FILL
XFILL_85_DFFSR_131 gnd vdd FILL
XFILL_1_DFFSR_235 gnd vdd FILL
XFILL_74_DFFSR_37 gnd vdd FILL
XFILL_12_OAI21X1_31 gnd vdd FILL
XFILL_9_4 gnd vdd FILL
XFILL_85_DFFSR_142 gnd vdd FILL
XFILL_74_DFFSR_48 gnd vdd FILL
XFILL_12_OAI21X1_42 gnd vdd FILL
XFILL_1_DFFSR_246 gnd vdd FILL
XFILL_85_DFFSR_153 gnd vdd FILL
XFILL_17_MUX2X1_5 gnd vdd FILL
XFILL_1_DFFSR_257 gnd vdd FILL
XFILL_74_DFFSR_59 gnd vdd FILL
XFILL_1_DFFSR_268 gnd vdd FILL
XFILL_85_DFFSR_164 gnd vdd FILL
XFILL_1_NOR2X1_170 gnd vdd FILL
XFILL_85_DFFSR_175 gnd vdd FILL
XFILL_17_CLKBUF1_4 gnd vdd FILL
XFILL_5_DFFSR_201 gnd vdd FILL
XFILL_85_DFFSR_186 gnd vdd FILL
XFILL_1_NOR2X1_181 gnd vdd FILL
XFILL_85_DFFSR_197 gnd vdd FILL
XFILL_5_DFFSR_212 gnd vdd FILL
XFILL_2_NAND3X1_1 gnd vdd FILL
XFILL_1_NOR2X1_192 gnd vdd FILL
XFILL_5_DFFSR_223 gnd vdd FILL
XFILL_58_5 gnd vdd FILL
XFILL_5_DFFSR_234 gnd vdd FILL
XFILL_5_DFFSR_245 gnd vdd FILL
XFILL_8_BUFX4_60 gnd vdd FILL
XFILL_43_DFFSR_14 gnd vdd FILL
XFILL_5_DFFSR_256 gnd vdd FILL
XFILL_5_DFFSR_267 gnd vdd FILL
XFILL_8_BUFX4_71 gnd vdd FILL
XFILL_43_DFFSR_25 gnd vdd FILL
XFILL_8_BUFX4_82 gnd vdd FILL
XFILL_43_DFFSR_36 gnd vdd FILL
XFILL_63_6_1 gnd vdd FILL
XFILL_9_DFFSR_200 gnd vdd FILL
XFILL_8_BUFX4_93 gnd vdd FILL
XFILL_43_DFFSR_47 gnd vdd FILL
XFILL_9_DFFSR_211 gnd vdd FILL
XFILL_43_DFFSR_58 gnd vdd FILL
XFILL_9_DFFSR_222 gnd vdd FILL
XFILL_43_DFFSR_69 gnd vdd FILL
XFILL_62_1_0 gnd vdd FILL
XFILL_9_DFFSR_233 gnd vdd FILL
XFILL_9_DFFSR_244 gnd vdd FILL
XFILL_83_DFFSR_13 gnd vdd FILL
XFILL_9_DFFSR_255 gnd vdd FILL
XFILL_10_NAND3X1_109 gnd vdd FILL
XFILL_83_DFFSR_24 gnd vdd FILL
XFILL_9_DFFSR_266 gnd vdd FILL
XFILL_83_DFFSR_35 gnd vdd FILL
XFILL_1_MUX2X1_110 gnd vdd FILL
XFILL_83_DFFSR_46 gnd vdd FILL
XFILL_1_MUX2X1_121 gnd vdd FILL
XFILL_12_DFFSR_13 gnd vdd FILL
XFILL_67_DFFSR_109 gnd vdd FILL
XFILL_83_DFFSR_57 gnd vdd FILL
XFILL_83_DFFSR_68 gnd vdd FILL
XFILL_12_DFFSR_24 gnd vdd FILL
XFILL_1_MUX2X1_132 gnd vdd FILL
XFILL_83_DFFSR_79 gnd vdd FILL
XFILL_12_DFFSR_35 gnd vdd FILL
XFILL_1_MUX2X1_143 gnd vdd FILL
XFILL_12_DFFSR_46 gnd vdd FILL
XFILL_1_MUX2X1_154 gnd vdd FILL
XFILL_1_MUX2X1_165 gnd vdd FILL
XFILL_12_DFFSR_57 gnd vdd FILL
XFILL_14_NAND3X1_18 gnd vdd FILL
XFILL_12_DFFSR_68 gnd vdd FILL
XFILL_14_NAND3X1_29 gnd vdd FILL
XFILL_1_MUX2X1_176 gnd vdd FILL
XFILL_12_DFFSR_79 gnd vdd FILL
XFILL_1_MUX2X1_187 gnd vdd FILL
XFILL_52_DFFSR_12 gnd vdd FILL
XFILL_34_CLKBUF1_18 gnd vdd FILL
XFILL_52_DFFSR_23 gnd vdd FILL
XFILL_21_DFFSR_210 gnd vdd FILL
XFILL_52_DFFSR_34 gnd vdd FILL
XFILL_11_NOR2X1_12 gnd vdd FILL
XFILL_34_CLKBUF1_29 gnd vdd FILL
XFILL_23_NOR3X1_9 gnd vdd FILL
XFILL_21_DFFSR_221 gnd vdd FILL
XFILL_2_AOI22X1_6 gnd vdd FILL
XFILL_52_DFFSR_45 gnd vdd FILL
XFILL_11_NOR2X1_23 gnd vdd FILL
XFILL_52_DFFSR_56 gnd vdd FILL
XFILL_14_OAI21X1_9 gnd vdd FILL
XFILL_21_DFFSR_232 gnd vdd FILL
XFILL_11_NOR2X1_34 gnd vdd FILL
XFILL_21_DFFSR_243 gnd vdd FILL
XFILL_52_DFFSR_67 gnd vdd FILL
XFILL_11_NOR2X1_45 gnd vdd FILL
XFILL_11_NOR2X1_56 gnd vdd FILL
XFILL_52_DFFSR_78 gnd vdd FILL
XFILL_21_DFFSR_254 gnd vdd FILL
XFILL_52_DFFSR_89 gnd vdd FILL
XFILL_21_DFFSR_265 gnd vdd FILL
XFILL_11_NOR2X1_67 gnd vdd FILL
XFILL_11_NOR2X1_78 gnd vdd FILL
XFILL_2_INVX1_205 gnd vdd FILL
XFILL_2_INVX1_216 gnd vdd FILL
XFILL_9_MUX2X1_4 gnd vdd FILL
XFILL_11_NOR2X1_89 gnd vdd FILL
XFILL_1_DFFSR_7 gnd vdd FILL
XFILL_25_DFFSR_220 gnd vdd FILL
XFILL_2_INVX1_227 gnd vdd FILL
XFILL_14_DFFSR_5 gnd vdd FILL
XFILL_6_AOI22X1_5 gnd vdd FILL
XFILL_25_DFFSR_231 gnd vdd FILL
XFILL_21_DFFSR_11 gnd vdd FILL
XFILL_23_10 gnd vdd FILL
XFILL_25_DFFSR_242 gnd vdd FILL
XFILL_71_DFFSR_6 gnd vdd FILL
XFILL_21_DFFSR_22 gnd vdd FILL
XFILL_25_DFFSR_253 gnd vdd FILL
XFILL_21_DFFSR_33 gnd vdd FILL
XFILL_25_DFFSR_264 gnd vdd FILL
XFILL_21_DFFSR_44 gnd vdd FILL
XFILL_25_DFFSR_275 gnd vdd FILL
XFILL_21_DFFSR_55 gnd vdd FILL
XFILL_6_INVX1_204 gnd vdd FILL
XFILL_6_INVX1_215 gnd vdd FILL
XFILL_21_DFFSR_66 gnd vdd FILL
XFILL_21_DFFSR_77 gnd vdd FILL
XFILL_6_INVX1_226 gnd vdd FILL
XFILL_52_DFFSR_120 gnd vdd FILL
XFILL_21_DFFSR_88 gnd vdd FILL
XFILL_52_DFFSR_131 gnd vdd FILL
XFILL_21_DFFSR_99 gnd vdd FILL
XFILL_29_DFFSR_230 gnd vdd FILL
XFILL_52_DFFSR_142 gnd vdd FILL
XFILL_29_DFFSR_241 gnd vdd FILL
XFILL_61_DFFSR_10 gnd vdd FILL
XFILL_61_DFFSR_21 gnd vdd FILL
XFILL_52_DFFSR_153 gnd vdd FILL
XFILL_29_DFFSR_252 gnd vdd FILL
XFILL_61_DFFSR_32 gnd vdd FILL
XFILL_61_DFFSR_43 gnd vdd FILL
XFILL_29_DFFSR_263 gnd vdd FILL
XFILL_52_DFFSR_164 gnd vdd FILL
XFILL_29_DFFSR_274 gnd vdd FILL
XFILL_52_DFFSR_175 gnd vdd FILL
XFILL_61_DFFSR_54 gnd vdd FILL
XFILL_52_DFFSR_186 gnd vdd FILL
XFILL_52_DFFSR_197 gnd vdd FILL
XFILL_61_DFFSR_65 gnd vdd FILL
XFILL_61_DFFSR_76 gnd vdd FILL
XFILL_61_DFFSR_87 gnd vdd FILL
XFILL_4_NAND3X1_13 gnd vdd FILL
XFILL_56_DFFSR_130 gnd vdd FILL
XFILL_61_DFFSR_98 gnd vdd FILL
XFILL_4_NAND3X1_24 gnd vdd FILL
XFILL_54_6_1 gnd vdd FILL
XFILL_4_NAND3X1_35 gnd vdd FILL
XFILL_56_DFFSR_141 gnd vdd FILL
XFILL_56_DFFSR_152 gnd vdd FILL
XFILL_4_NAND3X1_46 gnd vdd FILL
XFILL_4_DFFSR_12 gnd vdd FILL
XFILL_56_DFFSR_163 gnd vdd FILL
XFILL_4_NAND3X1_57 gnd vdd FILL
XFILL_53_1_0 gnd vdd FILL
XFILL_4_DFFSR_23 gnd vdd FILL
XFILL_8_NAND2X1_15 gnd vdd FILL
XFILL_56_DFFSR_174 gnd vdd FILL
XFILL_8_NAND2X1_26 gnd vdd FILL
XFILL_4_NAND3X1_68 gnd vdd FILL
XFILL_4_DFFSR_34 gnd vdd FILL
XFILL_4_NAND3X1_79 gnd vdd FILL
XFILL_4_DFFSR_45 gnd vdd FILL
XFILL_56_DFFSR_185 gnd vdd FILL
XFILL_36_DFFSR_9 gnd vdd FILL
XFILL_30_DFFSR_20 gnd vdd FILL
XFILL_8_NAND2X1_37 gnd vdd FILL
XFILL_56_DFFSR_196 gnd vdd FILL
XFILL_4_DFFSR_56 gnd vdd FILL
XFILL_8_NAND2X1_48 gnd vdd FILL
XFILL_30_DFFSR_31 gnd vdd FILL
XFILL_8_NAND2X1_59 gnd vdd FILL
XFILL_4_DFFSR_67 gnd vdd FILL
XFILL_30_DFFSR_42 gnd vdd FILL
XFILL_4_DFFSR_78 gnd vdd FILL
XFILL_30_DFFSR_53 gnd vdd FILL
XFILL_4_DFFSR_89 gnd vdd FILL
XFILL_30_DFFSR_64 gnd vdd FILL
XFILL_30_DFFSR_75 gnd vdd FILL
XFILL_30_DFFSR_86 gnd vdd FILL
XFILL_3_DFFSR_100 gnd vdd FILL
XFILL_30_DFFSR_97 gnd vdd FILL
XFILL_3_DFFSR_111 gnd vdd FILL
XFILL_34_DFFSR_109 gnd vdd FILL
XFILL_70_DFFSR_30 gnd vdd FILL
XFILL_3_DFFSR_122 gnd vdd FILL
XFILL_3_DFFSR_133 gnd vdd FILL
XFILL_18_MUX2X1_190 gnd vdd FILL
XFILL_70_DFFSR_41 gnd vdd FILL
XFILL_3_DFFSR_144 gnd vdd FILL
XFILL_70_DFFSR_52 gnd vdd FILL
XFILL_70_DFFSR_63 gnd vdd FILL
XFILL_3_DFFSR_155 gnd vdd FILL
XFILL_70_DFFSR_74 gnd vdd FILL
XFILL_3_DFFSR_166 gnd vdd FILL
XFILL_3_DFFSR_177 gnd vdd FILL
XFILL_70_DFFSR_85 gnd vdd FILL
XFILL_70_DFFSR_96 gnd vdd FILL
XFILL_3_DFFSR_188 gnd vdd FILL
XFILL_7_DFFSR_110 gnd vdd FILL
XFILL_3_DFFSR_199 gnd vdd FILL
XFILL_38_DFFSR_108 gnd vdd FILL
XFILL_7_DFFSR_121 gnd vdd FILL
XFILL_7_DFFSR_132 gnd vdd FILL
XFILL_11_MUX2X1_30 gnd vdd FILL
XFILL_38_DFFSR_119 gnd vdd FILL
XFILL_7_DFFSR_143 gnd vdd FILL
XFILL_11_MUX2X1_41 gnd vdd FILL
XFILL_7_DFFSR_154 gnd vdd FILL
XFILL_11_MUX2X1_52 gnd vdd FILL
XFILL_7_DFFSR_165 gnd vdd FILL
XFILL_11_MUX2X1_63 gnd vdd FILL
XFILL_10_NOR3X1_4 gnd vdd FILL
XDFFSR_190 INVX1_96/A DFFSR_90/CLK BUFX4_21/Y vdd MUX2X1_83/Y gnd vdd DFFSR
XFILL_11_MUX2X1_74 gnd vdd FILL
XFILL_7_DFFSR_176 gnd vdd FILL
XFILL_11_MUX2X1_85 gnd vdd FILL
XFILL_7_DFFSR_187 gnd vdd FILL
XFILL_11_MUX2X1_96 gnd vdd FILL
XFILL_7_DFFSR_198 gnd vdd FILL
XFILL_15_MUX2X1_40 gnd vdd FILL
XFILL_15_MUX2X1_51 gnd vdd FILL
XFILL_15_MUX2X1_62 gnd vdd FILL
XFILL_15_MUX2X1_73 gnd vdd FILL
XFILL_3_NOR3X1_11 gnd vdd FILL
XFILL_15_MUX2X1_84 gnd vdd FILL
XFILL_3_NOR3X1_22 gnd vdd FILL
XFILL_3_NOR3X1_33 gnd vdd FILL
XFILL_15_MUX2X1_95 gnd vdd FILL
XFILL_3_NOR3X1_44 gnd vdd FILL
XFILL_23_CLKBUF1_14 gnd vdd FILL
XFILL_23_CLKBUF1_25 gnd vdd FILL
XFILL_84_DFFSR_209 gnd vdd FILL
XFILL_23_CLKBUF1_36 gnd vdd FILL
XFILL_19_MUX2X1_50 gnd vdd FILL
XFILL_19_MUX2X1_61 gnd vdd FILL
XFILL_19_MUX2X1_72 gnd vdd FILL
XFILL_7_NOR3X1_10 gnd vdd FILL
XFILL_19_MUX2X1_83 gnd vdd FILL
XFILL_7_NOR3X1_21 gnd vdd FILL
XFILL_0_INVX1_104 gnd vdd FILL
XFILL_19_MUX2X1_94 gnd vdd FILL
XFILL_6_CLKBUF1_18 gnd vdd FILL
XFILL_7_NOR3X1_32 gnd vdd FILL
XFILL_6_CLKBUF1_29 gnd vdd FILL
XFILL_7_NOR3X1_43 gnd vdd FILL
XFILL_0_INVX1_115 gnd vdd FILL
XFILL_45_6_1 gnd vdd FILL
XFILL_0_INVX1_126 gnd vdd FILL
XFILL_1_AOI21X1_15 gnd vdd FILL
XFILL_0_INVX1_137 gnd vdd FILL
XFILL_23_DFFSR_130 gnd vdd FILL
XFILL_44_1_0 gnd vdd FILL
XFILL_1_AOI21X1_26 gnd vdd FILL
XFILL_0_INVX1_148 gnd vdd FILL
XFILL_23_DFFSR_141 gnd vdd FILL
XFILL_0_INVX1_159 gnd vdd FILL
XFILL_23_DFFSR_152 gnd vdd FILL
XFILL_1_AOI21X1_37 gnd vdd FILL
XFILL_23_DFFSR_163 gnd vdd FILL
XFILL_1_AOI21X1_48 gnd vdd FILL
XFILL_1_AOI21X1_59 gnd vdd FILL
XFILL_23_DFFSR_174 gnd vdd FILL
XFILL_11_OAI22X1_17 gnd vdd FILL
XFILL_4_INVX1_103 gnd vdd FILL
XFILL_4_INVX1_114 gnd vdd FILL
XFILL_11_OAI22X1_28 gnd vdd FILL
XFILL_23_DFFSR_185 gnd vdd FILL
XFILL_11_OAI22X1_39 gnd vdd FILL
XFILL_23_DFFSR_196 gnd vdd FILL
XFILL_4_INVX1_125 gnd vdd FILL
XFILL_4_NOR2X1_103 gnd vdd FILL
XFILL_4_NOR2X1_114 gnd vdd FILL
XFILL_4_INVX1_136 gnd vdd FILL
XFILL_4_INVX1_147 gnd vdd FILL
XFILL_15_OAI21X1_19 gnd vdd FILL
XFILL_4_NOR2X1_125 gnd vdd FILL
XFILL_27_DFFSR_140 gnd vdd FILL
XFILL_4_INVX1_158 gnd vdd FILL
XFILL_27_DFFSR_151 gnd vdd FILL
XFILL_4_NOR2X1_136 gnd vdd FILL
XFILL_27_DFFSR_162 gnd vdd FILL
XFILL_4_NOR2X1_147 gnd vdd FILL
XFILL_4_INVX1_169 gnd vdd FILL
XFILL_4_NOR2X1_158 gnd vdd FILL
XFILL_27_DFFSR_173 gnd vdd FILL
XFILL_4_NOR2X1_169 gnd vdd FILL
XFILL_27_DFFSR_184 gnd vdd FILL
XFILL_10_NAND3X1_60 gnd vdd FILL
XFILL_27_DFFSR_195 gnd vdd FILL
XFILL_10_NAND3X1_71 gnd vdd FILL
XFILL_2_NOR3X1_3 gnd vdd FILL
XFILL_10_NAND3X1_82 gnd vdd FILL
XFILL_11_INVX8_3 gnd vdd FILL
XFILL_10_NAND3X1_93 gnd vdd FILL
XFILL_23_NOR3X1_30 gnd vdd FILL
XFILL_23_NOR3X1_41 gnd vdd FILL
XFILL_21_MUX2X1_105 gnd vdd FILL
XFILL_23_NOR3X1_52 gnd vdd FILL
XFILL_21_MUX2X1_116 gnd vdd FILL
XFILL_21_MUX2X1_127 gnd vdd FILL
XFILL_73_DFFSR_230 gnd vdd FILL
XFILL_2_OAI22X1_9 gnd vdd FILL
XFILL_21_MUX2X1_138 gnd vdd FILL
XFILL_21_MUX2X1_149 gnd vdd FILL
XFILL_73_DFFSR_241 gnd vdd FILL
XFILL_73_DFFSR_252 gnd vdd FILL
XFILL_0_DFFSR_60 gnd vdd FILL
XFILL_73_DFFSR_263 gnd vdd FILL
XFILL_53_DFFSR_3 gnd vdd FILL
XFILL_73_DFFSR_274 gnd vdd FILL
XFILL_4_MUX2X1_109 gnd vdd FILL
XFILL_27_NOR3X1_40 gnd vdd FILL
XFILL_0_DFFSR_71 gnd vdd FILL
XFILL_0_DFFSR_82 gnd vdd FILL
XFILL_27_NOR3X1_51 gnd vdd FILL
XFILL_7_1 gnd vdd FILL
XFILL_0_DFFSR_93 gnd vdd FILL
XFILL_9_NOR2X1_203 gnd vdd FILL
XFILL_6_OAI22X1_8 gnd vdd FILL
XFILL_1_OAI22X1_12 gnd vdd FILL
XFILL_1_OAI22X1_23 gnd vdd FILL
XFILL_77_DFFSR_240 gnd vdd FILL
XFILL_63_3 gnd vdd FILL
XFILL_1_OAI22X1_34 gnd vdd FILL
XFILL_77_DFFSR_251 gnd vdd FILL
XFILL_77_DFFSR_262 gnd vdd FILL
XFILL_1_OAI22X1_45 gnd vdd FILL
XFILL_32_CLKBUF1_3 gnd vdd FILL
XFILL_5_OAI21X1_14 gnd vdd FILL
XFILL_77_DFFSR_273 gnd vdd FILL
XFILL_56_2 gnd vdd FILL
XFILL_5_OAI21X1_25 gnd vdd FILL
XFILL_5_OAI21X1_36 gnd vdd FILL
XFILL_51_DFFSR_209 gnd vdd FILL
XFILL_5_OAI21X1_47 gnd vdd FILL
XFILL_36_6_1 gnd vdd FILL
XFILL_35_1_0 gnd vdd FILL
XFILL_5_DFFSR_8 gnd vdd FILL
XFILL_55_DFFSR_208 gnd vdd FILL
XFILL_55_DFFSR_219 gnd vdd FILL
XFILL_18_DFFSR_6 gnd vdd FILL
XFILL_4_NAND2X1_90 gnd vdd FILL
XFILL_9_BUFX4_16 gnd vdd FILL
XFILL_75_DFFSR_7 gnd vdd FILL
XFILL_9_BUFX4_27 gnd vdd FILL
XFILL_9_BUFX4_38 gnd vdd FILL
XFILL_12_CLKBUF1_10 gnd vdd FILL
XFILL_9_BUFX4_49 gnd vdd FILL
XFILL_12_CLKBUF1_21 gnd vdd FILL
XFILL_82_DFFSR_108 gnd vdd FILL
XFILL_59_DFFSR_207 gnd vdd FILL
XFILL_12_CLKBUF1_32 gnd vdd FILL
XFILL_82_DFFSR_119 gnd vdd FILL
XFILL_59_DFFSR_218 gnd vdd FILL
XFILL_59_DFFSR_229 gnd vdd FILL
XFILL_86_DFFSR_107 gnd vdd FILL
XFILL_86_DFFSR_118 gnd vdd FILL
XFILL_86_DFFSR_129 gnd vdd FILL
XFILL_10_NOR2X1_150 gnd vdd FILL
XFILL_10_NOR2X1_161 gnd vdd FILL
XFILL_10_NOR2X1_172 gnd vdd FILL
XFILL_10_NOR2X1_183 gnd vdd FILL
XFILL_10_NOR2X1_194 gnd vdd FILL
XFILL_40_DFFSR_230 gnd vdd FILL
XFILL_40_DFFSR_241 gnd vdd FILL
XFILL_40_DFFSR_252 gnd vdd FILL
XNAND3X1_1 OAI21X1_1/A NAND3X1_1/B AND2X2_8/B gnd NAND3X1_1/Y vdd NAND3X1
XFILL_40_DFFSR_263 gnd vdd FILL
XFILL_40_DFFSR_274 gnd vdd FILL
XFILL_7_NAND3X1_9 gnd vdd FILL
XFILL_44_DFFSR_240 gnd vdd FILL
XFILL_13_BUFX4_10 gnd vdd FILL
XFILL_44_DFFSR_251 gnd vdd FILL
XFILL_44_DFFSR_262 gnd vdd FILL
XFILL_13_BUFX4_21 gnd vdd FILL
XFILL_44_DFFSR_273 gnd vdd FILL
XFILL_13_BUFX4_32 gnd vdd FILL
XFILL_27_6_1 gnd vdd FILL
XFILL_13_BUFX4_43 gnd vdd FILL
XFILL_2_6_1 gnd vdd FILL
XFILL_10_MUX2X1_101 gnd vdd FILL
XFILL_12_BUFX4_6 gnd vdd FILL
XFILL_10_MUX2X1_112 gnd vdd FILL
XFILL_13_BUFX4_54 gnd vdd FILL
XFILL_13_BUFX4_65 gnd vdd FILL
XFILL_26_1_0 gnd vdd FILL
XFILL_10_MUX2X1_123 gnd vdd FILL
XFILL_1_1_0 gnd vdd FILL
XFILL_71_DFFSR_140 gnd vdd FILL
XFILL_13_BUFX4_76 gnd vdd FILL
XFILL_10_MUX2X1_134 gnd vdd FILL
XFILL_10_MUX2X1_145 gnd vdd FILL
XFILL_71_DFFSR_151 gnd vdd FILL
XFILL_13_BUFX4_87 gnd vdd FILL
XFILL_71_DFFSR_162 gnd vdd FILL
XFILL_10_MUX2X1_156 gnd vdd FILL
XFILL_48_DFFSR_250 gnd vdd FILL
XFILL_13_BUFX4_98 gnd vdd FILL
XFILL_10_MUX2X1_167 gnd vdd FILL
XFILL_48_DFFSR_261 gnd vdd FILL
XFILL_48_DFFSR_272 gnd vdd FILL
XFILL_71_DFFSR_173 gnd vdd FILL
XFILL_71_DFFSR_184 gnd vdd FILL
XFILL_10_MUX2X1_178 gnd vdd FILL
XFILL_10_MUX2X1_189 gnd vdd FILL
XFILL_71_DFFSR_195 gnd vdd FILL
XFILL_22_DFFSR_208 gnd vdd FILL
XFILL_22_DFFSR_219 gnd vdd FILL
XFILL_11_OAI21X1_50 gnd vdd FILL
XFILL_75_DFFSR_150 gnd vdd FILL
XFILL_75_DFFSR_161 gnd vdd FILL
XFILL_75_DFFSR_172 gnd vdd FILL
XFILL_75_DFFSR_183 gnd vdd FILL
XFILL_75_DFFSR_194 gnd vdd FILL
XFILL_10_5_1 gnd vdd FILL
XFILL_26_DFFSR_207 gnd vdd FILL
XAOI22X1_6 AND2X2_4/Y NOR2X1_3/A DFFSR_275/Q INVX1_123/Y gnd AOI22X1_6/Y vdd AOI22X1
XFILL_26_DFFSR_218 gnd vdd FILL
XFILL_26_DFFSR_229 gnd vdd FILL
XFILL_7_INVX1_11 gnd vdd FILL
XFILL_79_DFFSR_160 gnd vdd FILL
XFILL_7_INVX1_22 gnd vdd FILL
XFILL_7_INVX1_33 gnd vdd FILL
XFILL_79_DFFSR_171 gnd vdd FILL
XINVX1_205 INVX1_205/A gnd INVX1_205/Y vdd INVX1
XFILL_7_INVX1_44 gnd vdd FILL
XFILL_79_DFFSR_182 gnd vdd FILL
XINVX1_216 DFFSR_69/Q gnd INVX1_216/Y vdd INVX1
XFILL_8_AND2X2_3 gnd vdd FILL
XFILL_53_DFFSR_107 gnd vdd FILL
XFILL_7_INVX1_55 gnd vdd FILL
XFILL_79_DFFSR_193 gnd vdd FILL
XINVX1_227 DFFSR_62/Q gnd INVX1_227/Y vdd INVX1
XFILL_7_INVX1_66 gnd vdd FILL
XFILL_7_INVX1_77 gnd vdd FILL
XFILL_53_DFFSR_118 gnd vdd FILL
XFILL_7_INVX1_88 gnd vdd FILL
XFILL_53_DFFSR_129 gnd vdd FILL
XFILL_71_DFFSR_19 gnd vdd FILL
XFILL_7_INVX1_99 gnd vdd FILL
XFILL_9_2_0 gnd vdd FILL
XFILL_14_MUX2X1_9 gnd vdd FILL
XFILL_57_DFFSR_106 gnd vdd FILL
XFILL_57_DFFSR_117 gnd vdd FILL
XFILL_0_MUX2X1_140 gnd vdd FILL
XFILL_57_DFFSR_128 gnd vdd FILL
XFILL_5_BUFX4_20 gnd vdd FILL
XFILL_57_DFFSR_139 gnd vdd FILL
XFILL_0_MUX2X1_151 gnd vdd FILL
XFILL_5_BUFX4_31 gnd vdd FILL
XFILL_0_MUX2X1_162 gnd vdd FILL
XFILL_13_NAND3X1_15 gnd vdd FILL
XNAND2X1_16 AND2X2_7/Y INVX2_1/A gnd NAND2X1_16/Y vdd NAND2X1
XFILL_0_MUX2X1_173 gnd vdd FILL
XNAND2X1_27 AND2X2_1/B NOR2X1_42/Y gnd NOR2X1_52/B vdd NAND2X1
XFILL_13_NAND3X1_26 gnd vdd FILL
XFILL_5_BUFX4_42 gnd vdd FILL
XFILL_13_NAND3X1_37 gnd vdd FILL
XFILL_0_MUX2X1_184 gnd vdd FILL
XFILL_5_BUFX4_53 gnd vdd FILL
XNAND2X1_38 NOR2X1_49/Y NOR2X1_48/Y gnd NOR3X1_3/B vdd NAND2X1
XNAND2X1_49 INVX1_100/A INVX1_125/Y gnd NAND3X1_65/A vdd NAND2X1
XFILL_5_BUFX4_64 gnd vdd FILL
XFILL_13_NAND3X1_48 gnd vdd FILL
XFILL_40_DFFSR_18 gnd vdd FILL
XFILL_13_NAND3X1_59 gnd vdd FILL
XFILL_5_BUFX4_75 gnd vdd FILL
XFILL_15_INVX8_4 gnd vdd FILL
XFILL_40_DFFSR_29 gnd vdd FILL
XFILL_33_CLKBUF1_15 gnd vdd FILL
XFILL_5_BUFX4_86 gnd vdd FILL
XFILL_33_CLKBUF1_26 gnd vdd FILL
XFILL_5_BUFX4_97 gnd vdd FILL
XFILL_33_CLKBUF1_37 gnd vdd FILL
XFILL_18_6_1 gnd vdd FILL
XFILL_11_DFFSR_240 gnd vdd FILL
XFILL_11_DFFSR_251 gnd vdd FILL
XFILL_11_DFFSR_262 gnd vdd FILL
XFILL_17_1_0 gnd vdd FILL
XFILL_4_DFFSR_109 gnd vdd FILL
XFILL_80_DFFSR_17 gnd vdd FILL
XFILL_11_DFFSR_273 gnd vdd FILL
XFILL_80_DFFSR_28 gnd vdd FILL
XFILL_80_DFFSR_39 gnd vdd FILL
XFILL_23_MUX2X1_7 gnd vdd FILL
XFILL_60_4_1 gnd vdd FILL
XFILL_28_6 gnd vdd FILL
XFILL_15_DFFSR_250 gnd vdd FILL
XFILL_15_DFFSR_261 gnd vdd FILL
XFILL_57_DFFSR_4 gnd vdd FILL
XFILL_8_DFFSR_108 gnd vdd FILL
XFILL_15_DFFSR_272 gnd vdd FILL
XFILL_8_DFFSR_119 gnd vdd FILL
XFILL_12_MUX2X1_17 gnd vdd FILL
XFILL_12_MUX2X1_28 gnd vdd FILL
XFILL_12_MUX2X1_39 gnd vdd FILL
XFILL_3_AOI21X1_4 gnd vdd FILL
XFILL_42_DFFSR_150 gnd vdd FILL
XFILL_42_DFFSR_161 gnd vdd FILL
XFILL_19_DFFSR_260 gnd vdd FILL
XFILL_19_DFFSR_271 gnd vdd FILL
XFILL_42_DFFSR_172 gnd vdd FILL
XFILL_42_DFFSR_183 gnd vdd FILL
XFILL_16_MUX2X1_16 gnd vdd FILL
XFILL_42_DFFSR_194 gnd vdd FILL
XFILL_16_MUX2X1_27 gnd vdd FILL
XFILL_3_NAND3X1_10 gnd vdd FILL
XFILL_16_MUX2X1_38 gnd vdd FILL
XFILL_3_NAND3X1_21 gnd vdd FILL
XFILL_7_AOI21X1_3 gnd vdd FILL
XFILL_16_MUX2X1_49 gnd vdd FILL
XFILL_6_MUX2X1_8 gnd vdd FILL
XFILL_3_NAND3X1_32 gnd vdd FILL
XFILL_3_NAND3X1_43 gnd vdd FILL
XNOR3X1_4 NOR3X1_4/A NOR3X1_4/B NOR3X1_6/C gnd NOR3X1_7/B vdd NOR3X1
XFILL_46_DFFSR_160 gnd vdd FILL
XFILL_3_NAND3X1_54 gnd vdd FILL
XFILL_7_NAND2X1_12 gnd vdd FILL
XFILL_46_DFFSR_171 gnd vdd FILL
XFILL_3_NAND3X1_65 gnd vdd FILL
XFILL_7_NAND2X1_23 gnd vdd FILL
XFILL_3_NAND3X1_76 gnd vdd FILL
XFILL_46_DFFSR_182 gnd vdd FILL
XFILL_7_NAND2X1_34 gnd vdd FILL
XFILL_20_DFFSR_107 gnd vdd FILL
XFILL_9_DFFSR_9 gnd vdd FILL
XFILL_3_NAND3X1_87 gnd vdd FILL
XFILL_46_DFFSR_193 gnd vdd FILL
XFILL_7_NAND2X1_45 gnd vdd FILL
XFILL_3_NAND3X1_98 gnd vdd FILL
XFILL_20_DFFSR_118 gnd vdd FILL
XFILL_7_NAND2X1_56 gnd vdd FILL
XFILL_20_DFFSR_129 gnd vdd FILL
XFILL_7_NAND2X1_67 gnd vdd FILL
XFILL_7_NAND2X1_78 gnd vdd FILL
XFILL_79_DFFSR_8 gnd vdd FILL
XFILL_7_NAND2X1_89 gnd vdd FILL
XFILL_8_NOR3X1_19 gnd vdd FILL
XFILL_24_DFFSR_106 gnd vdd FILL
XFILL_24_DFFSR_117 gnd vdd FILL
XFILL_24_DFFSR_128 gnd vdd FILL
XFILL_24_DFFSR_139 gnd vdd FILL
XFILL_10_AOI21X1_17 gnd vdd FILL
XFILL_10_AOI21X1_28 gnd vdd FILL
XFILL_10_AOI21X1_39 gnd vdd FILL
XFILL_28_DFFSR_105 gnd vdd FILL
XFILL_1_DFFSR_16 gnd vdd FILL
XFILL_28_DFFSR_116 gnd vdd FILL
XFILL_1_DFFSR_27 gnd vdd FILL
XFILL_1_DFFSR_38 gnd vdd FILL
XFILL_11_NOR2X1_4 gnd vdd FILL
XFILL_28_DFFSR_127 gnd vdd FILL
XFILL_1_DFFSR_49 gnd vdd FILL
XFILL_28_DFFSR_138 gnd vdd FILL
XFILL_28_DFFSR_149 gnd vdd FILL
XFILL_7_AOI22X1_10 gnd vdd FILL
XFILL_20_NOR3X1_18 gnd vdd FILL
XFILL_3_INVX1_70 gnd vdd FILL
XFILL_20_NOR3X1_29 gnd vdd FILL
XFILL_51_4_1 gnd vdd FILL
XFILL_3_INVX1_81 gnd vdd FILL
XFILL_3_INVX1_92 gnd vdd FILL
XFILL_70_DFFSR_207 gnd vdd FILL
XFILL_49_DFFSR_40 gnd vdd FILL
XFILL_70_DFFSR_218 gnd vdd FILL
XFILL_49_DFFSR_51 gnd vdd FILL
XFILL_70_DFFSR_229 gnd vdd FILL
XFILL_10_MUX2X1_2 gnd vdd FILL
XFILL_49_DFFSR_62 gnd vdd FILL
XFILL_49_DFFSR_73 gnd vdd FILL
XFILL_49_DFFSR_84 gnd vdd FILL
XFILL_24_NOR3X1_17 gnd vdd FILL
XFILL_49_DFFSR_95 gnd vdd FILL
XFILL_24_NOR3X1_28 gnd vdd FILL
XFILL_22_CLKBUF1_11 gnd vdd FILL
XFILL_24_NOR3X1_39 gnd vdd FILL
XFILL_22_CLKBUF1_22 gnd vdd FILL
XFILL_74_DFFSR_206 gnd vdd FILL
XFILL_74_DFFSR_217 gnd vdd FILL
XFILL_22_CLKBUF1_33 gnd vdd FILL
XFILL_74_DFFSR_228 gnd vdd FILL
XFILL_74_DFFSR_239 gnd vdd FILL
XFILL_28_NOR3X1_16 gnd vdd FILL
XFILL_3_BUFX4_9 gnd vdd FILL
XFILL_5_CLKBUF1_15 gnd vdd FILL
XFILL_28_NOR3X1_27 gnd vdd FILL
XFILL_1_BUFX4_90 gnd vdd FILL
XFILL_5_CLKBUF1_26 gnd vdd FILL
XFILL_18_DFFSR_50 gnd vdd FILL
XFILL_28_NOR3X1_38 gnd vdd FILL
XFILL_5_CLKBUF1_37 gnd vdd FILL
XFILL_18_DFFSR_61 gnd vdd FILL
XFILL_28_NOR3X1_49 gnd vdd FILL
XFILL_18_DFFSR_72 gnd vdd FILL
XFILL_18_DFFSR_83 gnd vdd FILL
XFILL_78_DFFSR_205 gnd vdd FILL
XFILL_0_AOI21X1_12 gnd vdd FILL
XFILL_78_DFFSR_216 gnd vdd FILL
XFILL_18_DFFSR_94 gnd vdd FILL
XOAI22X1_9 OAI22X1_9/A OAI22X1_9/B OAI22X1_9/C OAI22X1_9/D gnd OAI22X1_9/Y vdd OAI22X1
XFILL_0_AOI21X1_23 gnd vdd FILL
XFILL_0_AOI21X1_34 gnd vdd FILL
XFILL_78_DFFSR_227 gnd vdd FILL
XFILL_78_DFFSR_238 gnd vdd FILL
XFILL_13_DFFSR_160 gnd vdd FILL
XFILL_0_AOI21X1_45 gnd vdd FILL
XFILL_29_NOR3X1_2 gnd vdd FILL
XFILL_78_DFFSR_249 gnd vdd FILL
XFILL_10_OAI22X1_14 gnd vdd FILL
XFILL_0_AOI21X1_56 gnd vdd FILL
XFILL_13_DFFSR_171 gnd vdd FILL
XFILL_0_AOI21X1_67 gnd vdd FILL
XFILL_2_CLKBUF1_3 gnd vdd FILL
XFILL_0_AOI21X1_78 gnd vdd FILL
XFILL_10_OAI22X1_25 gnd vdd FILL
XFILL_13_DFFSR_182 gnd vdd FILL
XFILL_13_DFFSR_193 gnd vdd FILL
XFILL_10_OAI22X1_36 gnd vdd FILL
XFILL_58_DFFSR_60 gnd vdd FILL
XFILL_10_OAI22X1_47 gnd vdd FILL
XFILL_3_NOR2X1_100 gnd vdd FILL
XFILL_58_DFFSR_71 gnd vdd FILL
XFILL_58_DFFSR_82 gnd vdd FILL
XFILL_3_NOR2X1_111 gnd vdd FILL
XFILL_58_DFFSR_93 gnd vdd FILL
XFILL_14_OAI21X1_16 gnd vdd FILL
XFILL_3_NOR2X1_122 gnd vdd FILL
XFILL_14_OAI21X1_27 gnd vdd FILL
XFILL_3_NOR2X1_133 gnd vdd FILL
XFILL_14_OAI21X1_38 gnd vdd FILL
XFILL_59_5_1 gnd vdd FILL
XFILL_14_OAI21X1_49 gnd vdd FILL
XFILL_3_NOR2X1_144 gnd vdd FILL
XFILL_3_NOR2X1_3 gnd vdd FILL
XFILL_17_DFFSR_170 gnd vdd FILL
XFILL_3_NOR2X1_155 gnd vdd FILL
XFILL_6_CLKBUF1_2 gnd vdd FILL
XFILL_3_NOR2X1_166 gnd vdd FILL
XFILL_17_DFFSR_181 gnd vdd FILL
XFILL_58_0_0 gnd vdd FILL
XFILL_3_NOR2X1_177 gnd vdd FILL
XFILL_17_DFFSR_192 gnd vdd FILL
XFILL_3_NOR2X1_188 gnd vdd FILL
XFILL_3_NOR2X1_199 gnd vdd FILL
XFILL_27_DFFSR_70 gnd vdd FILL
XFILL_27_DFFSR_81 gnd vdd FILL
XFILL_27_DFFSR_92 gnd vdd FILL
XFILL_2_MUX2X1_1 gnd vdd FILL
XFILL_20_MUX2X1_102 gnd vdd FILL
XFILL_20_MUX2X1_113 gnd vdd FILL
XFILL_20_MUX2X1_124 gnd vdd FILL
XFILL_20_MUX2X1_135 gnd vdd FILL
XFILL_67_DFFSR_80 gnd vdd FILL
XFILL_20_MUX2X1_146 gnd vdd FILL
XFILL_42_4_1 gnd vdd FILL
XFILL_67_DFFSR_91 gnd vdd FILL
XFILL_20_MUX2X1_157 gnd vdd FILL
XFILL_63_DFFSR_260 gnd vdd FILL
XFILL_20_MUX2X1_168 gnd vdd FILL
XFILL_63_DFFSR_271 gnd vdd FILL
XFILL_3_MUX2X1_106 gnd vdd FILL
XFILL_3_MUX2X1_117 gnd vdd FILL
XFILL_20_MUX2X1_179 gnd vdd FILL
XFILL_39_DFFSR_1 gnd vdd FILL
XFILL_3_MUX2X1_128 gnd vdd FILL
XFILL_3_MUX2X1_139 gnd vdd FILL
XFILL_8_NOR2X1_200 gnd vdd FILL
XFILL_0_OAI22X1_20 gnd vdd FILL
XFILL_0_OAI22X1_31 gnd vdd FILL
XFILL_0_OAI22X1_42 gnd vdd FILL
XFILL_4_OAI21X1_11 gnd vdd FILL
XFILL_67_DFFSR_270 gnd vdd FILL
XFILL_4_OAI21X1_22 gnd vdd FILL
XFILL_0_NOR2X1_10 gnd vdd FILL
XFILL_41_DFFSR_206 gnd vdd FILL
XFILL_36_DFFSR_90 gnd vdd FILL
XFILL_0_NOR2X1_21 gnd vdd FILL
XFILL_4_OAI21X1_33 gnd vdd FILL
XFILL_41_DFFSR_217 gnd vdd FILL
XFILL_4_OAI21X1_44 gnd vdd FILL
XFILL_3_OAI21X1_7 gnd vdd FILL
XFILL_41_DFFSR_228 gnd vdd FILL
XFILL_0_NOR2X1_32 gnd vdd FILL
XFILL_0_NOR2X1_43 gnd vdd FILL
XFILL_0_NOR2X1_54 gnd vdd FILL
XFILL_41_DFFSR_239 gnd vdd FILL
XFILL_0_NOR2X1_65 gnd vdd FILL
XFILL_0_NOR2X1_76 gnd vdd FILL
XAOI21X1_80 NAND3X1_38/Y BUFX2_7/A AOI22X1_3/A gnd AOI22X1_3/C vdd AOI21X1
XFILL_0_NOR2X1_87 gnd vdd FILL
XFILL_0_NOR2X1_98 gnd vdd FILL
XFILL_45_DFFSR_205 gnd vdd FILL
XFILL_4_NOR2X1_20 gnd vdd FILL
XFILL_4_NOR2X1_31 gnd vdd FILL
XFILL_45_DFFSR_216 gnd vdd FILL
XFILL_23_DFFSR_7 gnd vdd FILL
XFILL_7_OAI21X1_6 gnd vdd FILL
XFILL_45_DFFSR_227 gnd vdd FILL
XFILL_4_NOR2X1_42 gnd vdd FILL
XFILL_80_DFFSR_8 gnd vdd FILL
XFILL_45_DFFSR_238 gnd vdd FILL
XFILL_4_NOR2X1_53 gnd vdd FILL
XFILL_45_DFFSR_249 gnd vdd FILL
XFILL_4_NOR2X1_64 gnd vdd FILL
XFILL_4_NOR2X1_75 gnd vdd FILL
XFILL_4_NOR2X1_86 gnd vdd FILL
XFILL_72_DFFSR_105 gnd vdd FILL
XFILL_4_NOR2X1_97 gnd vdd FILL
XFILL_72_DFFSR_116 gnd vdd FILL
XFILL_49_DFFSR_204 gnd vdd FILL
XFILL_49_DFFSR_215 gnd vdd FILL
XFILL_8_NOR2X1_30 gnd vdd FILL
XFILL_49_0_0 gnd vdd FILL
XFILL_72_DFFSR_127 gnd vdd FILL
XFILL_49_DFFSR_226 gnd vdd FILL
XFILL_11_CLKBUF1_40 gnd vdd FILL
XFILL_72_DFFSR_138 gnd vdd FILL
XFILL_8_NOR2X1_41 gnd vdd FILL
XFILL_49_DFFSR_237 gnd vdd FILL
XFILL_72_DFFSR_149 gnd vdd FILL
XFILL_8_NOR2X1_52 gnd vdd FILL
XFILL_12_OAI22X1_3 gnd vdd FILL
XFILL_49_DFFSR_248 gnd vdd FILL
XFILL_8_NOR2X1_63 gnd vdd FILL
XFILL_8_NOR2X1_74 gnd vdd FILL
XFILL_49_DFFSR_259 gnd vdd FILL
XFILL_8_NOR2X1_85 gnd vdd FILL
XFILL_76_DFFSR_104 gnd vdd FILL
XFILL_8_NOR2X1_96 gnd vdd FILL
XFILL_76_DFFSR_115 gnd vdd FILL
XFILL_76_DFFSR_126 gnd vdd FILL
XFILL_76_DFFSR_137 gnd vdd FILL
XFILL_16_OAI22X1_2 gnd vdd FILL
XFILL_76_DFFSR_148 gnd vdd FILL
XFILL_76_DFFSR_159 gnd vdd FILL
XFILL_33_4_1 gnd vdd FILL
XFILL_26_3 gnd vdd FILL
XFILL_30_DFFSR_260 gnd vdd FILL
XFILL_19_2 gnd vdd FILL
XFILL_30_DFFSR_271 gnd vdd FILL
XFILL_0_NAND2X1_9 gnd vdd FILL
XFILL_34_DFFSR_270 gnd vdd FILL
XFILL_4_NAND2X1_8 gnd vdd FILL
XFILL_0_MUX2X1_50 gnd vdd FILL
XFILL_0_MUX2X1_61 gnd vdd FILL
XFILL_0_MUX2X1_72 gnd vdd FILL
XFILL_0_MUX2X1_83 gnd vdd FILL
XFILL_13_AND2X2_8 gnd vdd FILL
XFILL_61_DFFSR_170 gnd vdd FILL
XFILL_0_MUX2X1_94 gnd vdd FILL
XFILL_61_DFFSR_181 gnd vdd FILL
XFILL_8_NAND2X1_7 gnd vdd FILL
XFILL_61_DFFSR_192 gnd vdd FILL
XFILL_12_DFFSR_205 gnd vdd FILL
XFILL_12_DFFSR_216 gnd vdd FILL
XFILL_12_DFFSR_227 gnd vdd FILL
XFILL_4_MUX2X1_60 gnd vdd FILL
XFILL_4_MUX2X1_71 gnd vdd FILL
XFILL_12_DFFSR_238 gnd vdd FILL
XFILL_4_MUX2X1_82 gnd vdd FILL
XFILL_12_DFFSR_249 gnd vdd FILL
XFILL_31_10 gnd vdd FILL
XFILL_4_MUX2X1_93 gnd vdd FILL
XFILL_65_DFFSR_180 gnd vdd FILL
XFILL_65_DFFSR_191 gnd vdd FILL
XFILL_10_BUFX4_14 gnd vdd FILL
XFILL_16_DFFSR_204 gnd vdd FILL
XFILL_13_NAND3X1_4 gnd vdd FILL
XFILL_16_DFFSR_215 gnd vdd FILL
XFILL_10_BUFX4_25 gnd vdd FILL
XFILL_16_DFFSR_226 gnd vdd FILL
XFILL_10_BUFX4_36 gnd vdd FILL
XFILL_10_BUFX4_47 gnd vdd FILL
XFILL_16_DFFSR_237 gnd vdd FILL
XFILL_8_MUX2X1_70 gnd vdd FILL
XFILL_8_MUX2X1_81 gnd vdd FILL
XFILL_10_BUFX4_58 gnd vdd FILL
XFILL_8_MUX2X1_92 gnd vdd FILL
XFILL_10_BUFX4_69 gnd vdd FILL
XFILL_16_DFFSR_248 gnd vdd FILL
XFILL_16_DFFSR_259 gnd vdd FILL
XFILL_69_DFFSR_190 gnd vdd FILL
XFILL_43_DFFSR_104 gnd vdd FILL
XFILL_43_DFFSR_115 gnd vdd FILL
XFILL_43_DFFSR_126 gnd vdd FILL
XFILL_43_DFFSR_137 gnd vdd FILL
XFILL_43_DFFSR_148 gnd vdd FILL
XFILL_43_DFFSR_159 gnd vdd FILL
XFILL_24_4_1 gnd vdd FILL
XFILL_47_DFFSR_103 gnd vdd FILL
XFILL_47_DFFSR_114 gnd vdd FILL
XFILL_40_DFFSR_1 gnd vdd FILL
XFILL_47_DFFSR_125 gnd vdd FILL
XFILL_47_DFFSR_136 gnd vdd FILL
XFILL_12_NAND3X1_12 gnd vdd FILL
XFILL_47_DFFSR_147 gnd vdd FILL
XFILL_47_DFFSR_158 gnd vdd FILL
XFILL_12_NAND3X1_23 gnd vdd FILL
XFILL_47_DFFSR_169 gnd vdd FILL
XFILL_12_NAND3X1_34 gnd vdd FILL
XFILL_20_MUX2X1_80 gnd vdd FILL
XFILL_12_NAND3X1_45 gnd vdd FILL
XFILL_20_MUX2X1_91 gnd vdd FILL
XFILL_4_INVX1_15 gnd vdd FILL
XFILL_12_NAND3X1_56 gnd vdd FILL
XFILL_4_INVX1_26 gnd vdd FILL
XFILL_32_CLKBUF1_12 gnd vdd FILL
XFILL_4_INVX1_37 gnd vdd FILL
XFILL_12_NAND3X1_67 gnd vdd FILL
XFILL_32_CLKBUF1_23 gnd vdd FILL
XFILL_12_NAND3X1_78 gnd vdd FILL
XFILL_32_CLKBUF1_34 gnd vdd FILL
XFILL_12_NAND3X1_89 gnd vdd FILL
XFILL_4_INVX1_48 gnd vdd FILL
XFILL_5_AND2X2_7 gnd vdd FILL
XFILL_4_INVX1_59 gnd vdd FILL
XFILL_3_BUFX2_6 gnd vdd FILL
XFILL_13_AOI22X1_9 gnd vdd FILL
XFILL_17_AOI22X1_8 gnd vdd FILL
XFILL_2_BUFX4_13 gnd vdd FILL
XFILL_62_DFFSR_5 gnd vdd FILL
XFILL_2_BUFX4_24 gnd vdd FILL
XFILL_2_BUFX4_35 gnd vdd FILL
XFILL_19_DFFSR_17 gnd vdd FILL
XFILL_2_BUFX4_46 gnd vdd FILL
XFILL_2_BUFX4_57 gnd vdd FILL
XFILL_19_DFFSR_28 gnd vdd FILL
XFILL_2_BUFX4_68 gnd vdd FILL
XFILL_7_5_1 gnd vdd FILL
XFILL_19_DFFSR_39 gnd vdd FILL
XFILL_2_BUFX4_79 gnd vdd FILL
XFILL_3_OAI22X1_19 gnd vdd FILL
XFILL_6_0_0 gnd vdd FILL
XFILL_32_DFFSR_180 gnd vdd FILL
XFILL_59_DFFSR_16 gnd vdd FILL
XFILL_32_DFFSR_191 gnd vdd FILL
XFILL_59_DFFSR_27 gnd vdd FILL
XFILL_59_DFFSR_38 gnd vdd FILL
XFILL_59_DFFSR_49 gnd vdd FILL
XFILL_2_NAND3X1_40 gnd vdd FILL
XFILL_2_NAND3X1_51 gnd vdd FILL
XFILL_2_NAND3X1_62 gnd vdd FILL
XFILL_6_NAND2X1_20 gnd vdd FILL
XFILL_2_NAND3X1_73 gnd vdd FILL
XFILL_6_NAND2X1_31 gnd vdd FILL
XFILL_10_DFFSR_104 gnd vdd FILL
XFILL_2_NAND3X1_84 gnd vdd FILL
XFILL_36_DFFSR_190 gnd vdd FILL
XFILL_6_NAND2X1_42 gnd vdd FILL
XFILL_2_NAND3X1_95 gnd vdd FILL
XFILL_10_DFFSR_115 gnd vdd FILL
XFILL_27_DFFSR_8 gnd vdd FILL
XFILL_6_NAND2X1_53 gnd vdd FILL
XFILL_15_4_1 gnd vdd FILL
XFILL_10_DFFSR_126 gnd vdd FILL
XFILL_6_NAND2X1_64 gnd vdd FILL
XFILL_84_DFFSR_9 gnd vdd FILL
XFILL_10_DFFSR_137 gnd vdd FILL
XFILL_6_NAND2X1_75 gnd vdd FILL
XMUX2X1_2 MUX2X1_2/A MUX2X1_2/B MUX2X1_2/S gnd MUX2X1_2/Y vdd MUX2X1
XFILL_10_DFFSR_148 gnd vdd FILL
XFILL_6_NAND2X1_86 gnd vdd FILL
XFILL_28_DFFSR_15 gnd vdd FILL
XFILL_28_DFFSR_26 gnd vdd FILL
XFILL_10_DFFSR_159 gnd vdd FILL
XFILL_28_DFFSR_37 gnd vdd FILL
XFILL_28_DFFSR_48 gnd vdd FILL
XFILL_14_DFFSR_103 gnd vdd FILL
XFILL_28_DFFSR_59 gnd vdd FILL
XFILL_14_DFFSR_114 gnd vdd FILL
XFILL_14_CLKBUF1_17 gnd vdd FILL
XFILL_14_CLKBUF1_28 gnd vdd FILL
XFILL_14_DFFSR_125 gnd vdd FILL
XFILL_14_DFFSR_136 gnd vdd FILL
XFILL_14_CLKBUF1_39 gnd vdd FILL
XFILL_68_DFFSR_14 gnd vdd FILL
XFILL_14_DFFSR_147 gnd vdd FILL
XFILL_14_DFFSR_158 gnd vdd FILL
XFILL_68_DFFSR_25 gnd vdd FILL
XFILL_68_DFFSR_36 gnd vdd FILL
XFILL_14_DFFSR_169 gnd vdd FILL
XFILL_68_DFFSR_47 gnd vdd FILL
XFILL_68_DFFSR_58 gnd vdd FILL
XFILL_18_DFFSR_102 gnd vdd FILL
XFILL_68_DFFSR_69 gnd vdd FILL
XFILL_18_DFFSR_113 gnd vdd FILL
XFILL_18_DFFSR_124 gnd vdd FILL
XFILL_1_INVX1_4 gnd vdd FILL
XFILL_18_DFFSR_135 gnd vdd FILL
XFILL_18_DFFSR_146 gnd vdd FILL
XFILL_18_DFFSR_157 gnd vdd FILL
XCLKBUF1_3 BUFX4_95/Y gnd DFFSR_4/CLK vdd CLKBUF1
XFILL_18_DFFSR_168 gnd vdd FILL
XFILL_18_DFFSR_179 gnd vdd FILL
XFILL_37_DFFSR_13 gnd vdd FILL
XFILL_10_NOR3X1_15 gnd vdd FILL
XFILL_10_NOR3X1_26 gnd vdd FILL
XFILL_37_DFFSR_24 gnd vdd FILL
XFILL_10_NOR3X1_37 gnd vdd FILL
XFILL_37_DFFSR_35 gnd vdd FILL
XFILL_37_DFFSR_46 gnd vdd FILL
XFILL_10_NOR3X1_48 gnd vdd FILL
XFILL_60_DFFSR_204 gnd vdd FILL
XFILL_60_DFFSR_215 gnd vdd FILL
XFILL_37_DFFSR_57 gnd vdd FILL
XFILL_37_DFFSR_68 gnd vdd FILL
XFILL_60_DFFSR_226 gnd vdd FILL
XFILL_60_DFFSR_237 gnd vdd FILL
XFILL_37_DFFSR_79 gnd vdd FILL
XFILL_60_DFFSR_248 gnd vdd FILL
XFILL_14_NOR3X1_14 gnd vdd FILL
XFILL_77_DFFSR_12 gnd vdd FILL
XFILL_60_DFFSR_259 gnd vdd FILL
XFILL_77_DFFSR_23 gnd vdd FILL
XFILL_14_NOR3X1_25 gnd vdd FILL
XFILL_14_NOR3X1_36 gnd vdd FILL
XFILL_14_NOR3X1_47 gnd vdd FILL
XFILL_77_DFFSR_34 gnd vdd FILL
XFILL_21_CLKBUF1_30 gnd vdd FILL
XFILL_64_DFFSR_203 gnd vdd FILL
XFILL_77_DFFSR_45 gnd vdd FILL
XFILL_77_DFFSR_56 gnd vdd FILL
XFILL_64_DFFSR_214 gnd vdd FILL
XFILL_21_CLKBUF1_41 gnd vdd FILL
XFILL_77_DFFSR_67 gnd vdd FILL
XFILL_64_DFFSR_225 gnd vdd FILL
XFILL_77_DFFSR_78 gnd vdd FILL
XFILL_64_DFFSR_236 gnd vdd FILL
XFILL_7_BUFX4_105 gnd vdd FILL
XFILL_65_3_1 gnd vdd FILL
XFILL_77_DFFSR_89 gnd vdd FILL
XFILL_64_DFFSR_247 gnd vdd FILL
XFILL_4_CLKBUF1_12 gnd vdd FILL
XFILL_18_NOR3X1_13 gnd vdd FILL
XFILL_64_DFFSR_258 gnd vdd FILL
XFILL_0_INVX1_30 gnd vdd FILL
XFILL_64_DFFSR_269 gnd vdd FILL
XFILL_4_CLKBUF1_23 gnd vdd FILL
XFILL_18_NOR3X1_24 gnd vdd FILL
XFILL_0_INVX1_41 gnd vdd FILL
XFILL_4_CLKBUF1_34 gnd vdd FILL
XFILL_18_NOR3X1_35 gnd vdd FILL
XFILL_0_INVX1_52 gnd vdd FILL
XFILL_68_DFFSR_202 gnd vdd FILL
XFILL_18_NOR3X1_46 gnd vdd FILL
XNOR2X1_201 DFFSR_8/Q NOR2X1_202/B gnd NOR2X1_201/Y vdd NOR2X1
XFILL_0_INVX1_63 gnd vdd FILL
XFILL_12_MUX2X1_108 gnd vdd FILL
XFILL_12_MUX2X1_119 gnd vdd FILL
XFILL_68_DFFSR_213 gnd vdd FILL
XFILL_46_DFFSR_11 gnd vdd FILL
XFILL_0_INVX1_74 gnd vdd FILL
XFILL_0_INVX1_85 gnd vdd FILL
XFILL_46_DFFSR_22 gnd vdd FILL
XFILL_68_DFFSR_224 gnd vdd FILL
XFILL_68_DFFSR_235 gnd vdd FILL
XFILL_0_INVX1_96 gnd vdd FILL
XFILL_46_DFFSR_33 gnd vdd FILL
XFILL_17_NOR3X1_8 gnd vdd FILL
XFILL_68_DFFSR_246 gnd vdd FILL
XFILL_31_1 gnd vdd FILL
XFILL_46_DFFSR_44 gnd vdd FILL
XFILL_46_DFFSR_55 gnd vdd FILL
XFILL_68_DFFSR_257 gnd vdd FILL
XFILL_68_DFFSR_268 gnd vdd FILL
XFILL_46_DFFSR_66 gnd vdd FILL
XFILL_46_DFFSR_77 gnd vdd FILL
XFILL_23_CLKBUF1_9 gnd vdd FILL
XFILL_46_DFFSR_88 gnd vdd FILL
XFILL_1_NOR2X1_19 gnd vdd FILL
XFILL_13_OAI21X1_13 gnd vdd FILL
XFILL_46_DFFSR_99 gnd vdd FILL
XFILL_86_DFFSR_10 gnd vdd FILL
XFILL_86_DFFSR_21 gnd vdd FILL
XFILL_13_OAI21X1_24 gnd vdd FILL
XFILL_2_NOR2X1_130 gnd vdd FILL
XFILL_13_OAI21X1_35 gnd vdd FILL
XFILL_86_DFFSR_32 gnd vdd FILL
XFILL_86_DFFSR_43 gnd vdd FILL
XFILL_2_NOR2X1_141 gnd vdd FILL
XFILL_13_OAI21X1_46 gnd vdd FILL
XFILL_2_NOR2X1_152 gnd vdd FILL
XFILL_15_DFFSR_10 gnd vdd FILL
XFILL_86_DFFSR_54 gnd vdd FILL
XFILL_2_NOR2X1_163 gnd vdd FILL
XFILL_15_DFFSR_21 gnd vdd FILL
XFILL_2_NOR2X1_174 gnd vdd FILL
XFILL_86_DFFSR_65 gnd vdd FILL
XFILL_86_DFFSR_76 gnd vdd FILL
XFILL_27_CLKBUF1_8 gnd vdd FILL
XFILL_15_DFFSR_32 gnd vdd FILL
XFILL_2_NOR2X1_185 gnd vdd FILL
XFILL_15_DFFSR_43 gnd vdd FILL
XFILL_86_DFFSR_87 gnd vdd FILL
XFILL_5_NOR2X1_18 gnd vdd FILL
XFILL_86_DFFSR_98 gnd vdd FILL
XFILL_2_NOR2X1_196 gnd vdd FILL
XFILL_5_NOR2X1_29 gnd vdd FILL
XFILL_15_DFFSR_54 gnd vdd FILL
XFILL_26_10 gnd vdd FILL
XFILL_15_DFFSR_65 gnd vdd FILL
XFILL_15_DFFSR_76 gnd vdd FILL
XFILL_15_DFFSR_87 gnd vdd FILL
XFILL_15_DFFSR_98 gnd vdd FILL
XFILL_55_DFFSR_20 gnd vdd FILL
XFILL_55_DFFSR_31 gnd vdd FILL
XFILL_26_NOR3X1_6 gnd vdd FILL
XFILL_55_DFFSR_42 gnd vdd FILL
XFILL_55_DFFSR_53 gnd vdd FILL
XFILL_9_NOR2X1_17 gnd vdd FILL
XFILL_9_NOR2X1_28 gnd vdd FILL
XFILL_9_NOR2X1_39 gnd vdd FILL
XFILL_55_DFFSR_64 gnd vdd FILL
XFILL_55_DFFSR_75 gnd vdd FILL
XFILL_55_DFFSR_86 gnd vdd FILL
XFILL_55_DFFSR_97 gnd vdd FILL
XFILL_2_MUX2X1_103 gnd vdd FILL
XFILL_2_MUX2X1_114 gnd vdd FILL
XFILL_0_NOR2X1_7 gnd vdd FILL
XFILL_2_MUX2X1_125 gnd vdd FILL
XFILL_44_DFFSR_2 gnd vdd FILL
XFILL_2_MUX2X1_136 gnd vdd FILL
XFILL_2_MUX2X1_147 gnd vdd FILL
XFILL_24_DFFSR_30 gnd vdd FILL
XFILL_2_MUX2X1_158 gnd vdd FILL
XFILL_24_DFFSR_41 gnd vdd FILL
XFILL_2_MUX2X1_169 gnd vdd FILL
XFILL_24_DFFSR_52 gnd vdd FILL
XFILL_24_DFFSR_63 gnd vdd FILL
XFILL_24_DFFSR_74 gnd vdd FILL
XFILL_24_DFFSR_85 gnd vdd FILL
XFILL_80_DFFSR_190 gnd vdd FILL
XFILL_24_DFFSR_96 gnd vdd FILL
XFILL_56_3_1 gnd vdd FILL
XFILL_3_OAI21X1_30 gnd vdd FILL
XFILL_31_DFFSR_203 gnd vdd FILL
XFILL_9_NOR3X1_7 gnd vdd FILL
XFILL_3_OAI21X1_41 gnd vdd FILL
XFILL_31_DFFSR_214 gnd vdd FILL
XFILL_31_DFFSR_225 gnd vdd FILL
XFILL_7_BUFX2_7 gnd vdd FILL
XFILL_64_DFFSR_40 gnd vdd FILL
XFILL_31_DFFSR_236 gnd vdd FILL
XFILL_64_DFFSR_51 gnd vdd FILL
XFILL_31_DFFSR_247 gnd vdd FILL
XFILL_64_DFFSR_62 gnd vdd FILL
XFILL_0_DFFSR_260 gnd vdd FILL
XFILL_0_DFFSR_271 gnd vdd FILL
XFILL_64_DFFSR_73 gnd vdd FILL
XFILL_31_DFFSR_258 gnd vdd FILL
XFILL_31_DFFSR_269 gnd vdd FILL
XFILL_64_DFFSR_84 gnd vdd FILL
XFILL_64_DFFSR_95 gnd vdd FILL
XFILL_35_DFFSR_202 gnd vdd FILL
XFILL_35_DFFSR_213 gnd vdd FILL
XFILL_35_DFFSR_224 gnd vdd FILL
XFILL_35_DFFSR_235 gnd vdd FILL
XFILL_7_DFFSR_20 gnd vdd FILL
XFILL_7_DFFSR_31 gnd vdd FILL
XFILL_35_DFFSR_246 gnd vdd FILL
XFILL_7_DFFSR_42 gnd vdd FILL
XFILL_4_DFFSR_270 gnd vdd FILL
XFILL_66_DFFSR_6 gnd vdd FILL
XFILL_7_DFFSR_53 gnd vdd FILL
XFILL_35_DFFSR_257 gnd vdd FILL
XFILL_35_DFFSR_268 gnd vdd FILL
XFILL_1_MUX2X1_15 gnd vdd FILL
XFILL_7_DFFSR_64 gnd vdd FILL
XFILL_40_7_2 gnd vdd FILL
XFILL_1_MUX2X1_26 gnd vdd FILL
XFILL_39_DFFSR_201 gnd vdd FILL
XFILL_62_DFFSR_102 gnd vdd FILL
XFILL_7_DFFSR_75 gnd vdd FILL
XFILL_33_DFFSR_50 gnd vdd FILL
XFILL_7_DFFSR_86 gnd vdd FILL
XFILL_1_MUX2X1_37 gnd vdd FILL
XFILL_62_DFFSR_113 gnd vdd FILL
XFILL_33_DFFSR_61 gnd vdd FILL
XFILL_62_DFFSR_124 gnd vdd FILL
XFILL_39_DFFSR_212 gnd vdd FILL
XFILL_1_MUX2X1_48 gnd vdd FILL
XFILL_33_DFFSR_72 gnd vdd FILL
XFILL_7_DFFSR_97 gnd vdd FILL
XFILL_33_DFFSR_83 gnd vdd FILL
XFILL_1_MUX2X1_59 gnd vdd FILL
XFILL_39_DFFSR_223 gnd vdd FILL
XFILL_39_DFFSR_234 gnd vdd FILL
XFILL_62_DFFSR_135 gnd vdd FILL
XFILL_62_DFFSR_146 gnd vdd FILL
XFILL_39_DFFSR_245 gnd vdd FILL
XFILL_33_DFFSR_94 gnd vdd FILL
XFILL_62_DFFSR_157 gnd vdd FILL
XFILL_39_DFFSR_256 gnd vdd FILL
XFILL_62_DFFSR_168 gnd vdd FILL
XFILL_39_DFFSR_267 gnd vdd FILL
XFILL_5_MUX2X1_14 gnd vdd FILL
XFILL_62_DFFSR_179 gnd vdd FILL
XFILL_5_MUX2X1_25 gnd vdd FILL
XFILL_66_DFFSR_101 gnd vdd FILL
XFILL_73_DFFSR_60 gnd vdd FILL
XFILL_5_MUX2X1_36 gnd vdd FILL
XFILL_66_DFFSR_112 gnd vdd FILL
XFILL_5_NAND3X1_17 gnd vdd FILL
XFILL_5_MUX2X1_47 gnd vdd FILL
XFILL_73_DFFSR_71 gnd vdd FILL
XFILL_66_DFFSR_123 gnd vdd FILL
XFILL_73_DFFSR_82 gnd vdd FILL
XFILL_66_DFFSR_134 gnd vdd FILL
XFILL_5_MUX2X1_58 gnd vdd FILL
XFILL_5_MUX2X1_69 gnd vdd FILL
XFILL_73_DFFSR_93 gnd vdd FILL
XFILL_5_NAND3X1_28 gnd vdd FILL
XFILL_66_DFFSR_145 gnd vdd FILL
XFILL_5_NAND3X1_39 gnd vdd FILL
XFILL_66_DFFSR_156 gnd vdd FILL
XFILL_66_DFFSR_167 gnd vdd FILL
XFILL_66_DFFSR_178 gnd vdd FILL
XFILL_9_MUX2X1_13 gnd vdd FILL
XFILL_9_NAND2X1_19 gnd vdd FILL
XFILL_6_BUFX4_1 gnd vdd FILL
XFILL_9_MUX2X1_24 gnd vdd FILL
XFILL_9_MUX2X1_35 gnd vdd FILL
XFILL_66_DFFSR_189 gnd vdd FILL
XFILL_9_MUX2X1_46 gnd vdd FILL
XFILL_13_NOR3X1_1 gnd vdd FILL
XFILL_9_MUX2X1_57 gnd vdd FILL
XFILL_9_MUX2X1_68 gnd vdd FILL
XFILL_9_MUX2X1_79 gnd vdd FILL
XFILL_13_OAI21X1_1 gnd vdd FILL
XFILL_42_DFFSR_70 gnd vdd FILL
XFILL_19_MUX2X1_150 gnd vdd FILL
XFILL_42_DFFSR_81 gnd vdd FILL
XFILL_19_MUX2X1_161 gnd vdd FILL
XFILL_42_DFFSR_92 gnd vdd FILL
XFILL_10_NOR2X1_70 gnd vdd FILL
XFILL_10_NOR2X1_81 gnd vdd FILL
XFILL_19_MUX2X1_172 gnd vdd FILL
XBUFX4_14 BUFX4_3/Y gnd DFFSR_2/R vdd BUFX4
XBUFX4_25 BUFX4_47/A gnd DFFSR_91/R vdd BUFX4
XFILL_19_MUX2X1_183 gnd vdd FILL
XFILL_10_NOR2X1_92 gnd vdd FILL
XFILL_19_MUX2X1_194 gnd vdd FILL
XBUFX4_36 BUFX4_62/Y gnd DFFSR_82/R vdd BUFX4
XBUFX4_47 BUFX4_47/A gnd DFFSR_93/R vdd BUFX4
XBUFX4_58 BUFX4_60/A gnd BUFX4_58/Y vdd BUFX4
XBUFX4_69 INVX8_1/Y gnd MUX2X1_1/A vdd BUFX4
XFILL_47_3_1 gnd vdd FILL
XFILL_82_DFFSR_80 gnd vdd FILL
XFILL_82_DFFSR_91 gnd vdd FILL
XFILL_21_MUX2X1_12 gnd vdd FILL
XFILL_21_MUX2X1_23 gnd vdd FILL
XFILL_5_INVX1_5 gnd vdd FILL
XFILL_11_DFFSR_80 gnd vdd FILL
XFILL_21_MUX2X1_34 gnd vdd FILL
XFILL_11_DFFSR_91 gnd vdd FILL
XFILL_21_MUX2X1_45 gnd vdd FILL
XFILL_21_MUX2X1_56 gnd vdd FILL
XFILL_21_MUX2X1_67 gnd vdd FILL
XFILL_21_MUX2X1_78 gnd vdd FILL
XFILL_21_MUX2X1_89 gnd vdd FILL
XFILL_51_DFFSR_90 gnd vdd FILL
XFILL_31_7_2 gnd vdd FILL
XFILL_30_2_1 gnd vdd FILL
XFILL_24_CLKBUF1_18 gnd vdd FILL
XFILL_24_CLKBUF1_29 gnd vdd FILL
XFILL_6_INVX4_1 gnd vdd FILL
XFILL_33_DFFSR_101 gnd vdd FILL
XFILL_10_NAND2X1_3 gnd vdd FILL
XFILL_33_DFFSR_112 gnd vdd FILL
XFILL_33_DFFSR_123 gnd vdd FILL
XFILL_2_AOI21X1_19 gnd vdd FILL
XFILL_33_DFFSR_134 gnd vdd FILL
XFILL_33_DFFSR_145 gnd vdd FILL
XFILL_33_DFFSR_156 gnd vdd FILL
XFILL_2_DFFSR_180 gnd vdd FILL
XFILL_33_DFFSR_167 gnd vdd FILL
XFILL_33_DFFSR_178 gnd vdd FILL
XFILL_2_DFFSR_191 gnd vdd FILL
XFILL_37_DFFSR_100 gnd vdd FILL
XFILL_33_DFFSR_189 gnd vdd FILL
XFILL_37_DFFSR_111 gnd vdd FILL
XFILL_5_NOR2X1_107 gnd vdd FILL
XFILL_37_DFFSR_122 gnd vdd FILL
XFILL_5_NOR2X1_118 gnd vdd FILL
XFILL_37_DFFSR_133 gnd vdd FILL
XFILL_5_NOR2X1_129 gnd vdd FILL
XFILL_37_DFFSR_144 gnd vdd FILL
XFILL_11_NAND3X1_20 gnd vdd FILL
XFILL_37_DFFSR_155 gnd vdd FILL
XFILL_11_NAND3X1_31 gnd vdd FILL
XFILL_37_DFFSR_166 gnd vdd FILL
XFILL_37_DFFSR_177 gnd vdd FILL
XFILL_6_DFFSR_190 gnd vdd FILL
XFILL_11_NAND3X1_42 gnd vdd FILL
XFILL_11_NAND3X1_53 gnd vdd FILL
XFILL_37_DFFSR_188 gnd vdd FILL
XFILL_3_DFFSR_90 gnd vdd FILL
XFILL_11_NAND3X1_64 gnd vdd FILL
XFILL_37_DFFSR_199 gnd vdd FILL
XFILL_31_CLKBUF1_20 gnd vdd FILL
XFILL_11_NAND3X1_75 gnd vdd FILL
XFILL_11_NAND3X1_86 gnd vdd FILL
XFILL_38_3_1 gnd vdd FILL
XFILL_31_CLKBUF1_31 gnd vdd FILL
XFILL_11_NAND3X1_97 gnd vdd FILL
XFILL_31_CLKBUF1_42 gnd vdd FILL
XFILL_83_DFFSR_201 gnd vdd FILL
XFILL_22_MUX2X1_109 gnd vdd FILL
XFILL_83_DFFSR_212 gnd vdd FILL
XFILL_10_DFFSR_5 gnd vdd FILL
XFILL_83_DFFSR_223 gnd vdd FILL
XFILL_83_DFFSR_234 gnd vdd FILL
XFILL_10_AOI21X1_8 gnd vdd FILL
XFILL_83_DFFSR_245 gnd vdd FILL
XFILL_83_DFFSR_256 gnd vdd FILL
XFILL_83_DFFSR_267 gnd vdd FILL
XFILL_22_7_2 gnd vdd FILL
XFILL_48_DFFSR_3 gnd vdd FILL
XFILL_87_DFFSR_200 gnd vdd FILL
XFILL_1_INVX1_19 gnd vdd FILL
XFILL_21_2_1 gnd vdd FILL
XFILL_87_DFFSR_211 gnd vdd FILL
XFILL_87_DFFSR_222 gnd vdd FILL
XFILL_14_AOI21X1_7 gnd vdd FILL
XFILL_87_DFFSR_233 gnd vdd FILL
XFILL_2_OAI22X1_16 gnd vdd FILL
XFILL_87_DFFSR_244 gnd vdd FILL
XFILL_2_OAI22X1_27 gnd vdd FILL
XFILL_87_DFFSR_255 gnd vdd FILL
XFILL_2_OAI22X1_38 gnd vdd FILL
XFILL_2_OAI22X1_49 gnd vdd FILL
XFILL_87_DFFSR_266 gnd vdd FILL
XFILL_6_OAI21X1_18 gnd vdd FILL
XFILL_6_OAI21X1_29 gnd vdd FILL
XFILL_3_INVX1_150 gnd vdd FILL
XFILL_3_INVX1_161 gnd vdd FILL
XFILL_3_INVX1_172 gnd vdd FILL
XFILL_3_INVX1_183 gnd vdd FILL
XFILL_1_NAND3X1_70 gnd vdd FILL
XFILL_3_INVX1_194 gnd vdd FILL
XFILL_1_NAND3X1_81 gnd vdd FILL
XFILL_32_DFFSR_9 gnd vdd FILL
XFILL_1_NAND3X1_92 gnd vdd FILL
XFILL_5_NAND2X1_50 gnd vdd FILL
XFILL_5_NAND2X1_61 gnd vdd FILL
XFILL_5_NAND2X1_72 gnd vdd FILL
XFILL_7_INVX1_160 gnd vdd FILL
XFILL_5_NAND2X1_83 gnd vdd FILL
XFILL_7_INVX1_171 gnd vdd FILL
XFILL_5_NAND2X1_94 gnd vdd FILL
XFILL_7_INVX1_182 gnd vdd FILL
XFILL_7_INVX1_193 gnd vdd FILL
XFILL_13_CLKBUF1_14 gnd vdd FILL
XFILL_13_CLKBUF1_25 gnd vdd FILL
XFILL_13_CLKBUF1_36 gnd vdd FILL
XFILL_1_OAI22X1_1 gnd vdd FILL
XFILL_29_3_1 gnd vdd FILL
XFILL_4_3_1 gnd vdd FILL
XFILL_11_NOR2X1_110 gnd vdd FILL
XFILL_11_NOR2X1_121 gnd vdd FILL
XFILL_11_NOR2X1_132 gnd vdd FILL
XFILL_25_DFFSR_19 gnd vdd FILL
XFILL_11_NOR2X1_143 gnd vdd FILL
XFILL_11_NOR2X1_154 gnd vdd FILL
XFILL_11_NOR2X1_165 gnd vdd FILL
XFILL_50_DFFSR_201 gnd vdd FILL
XFILL_11_NOR2X1_176 gnd vdd FILL
XFILL_11_NOR2X1_187 gnd vdd FILL
XFILL_50_DFFSR_212 gnd vdd FILL
XFILL_11_NOR2X1_198 gnd vdd FILL
XFILL_50_DFFSR_223 gnd vdd FILL
XFILL_50_DFFSR_234 gnd vdd FILL
XFILL_13_7_2 gnd vdd FILL
XFILL_9_AOI21X1_50 gnd vdd FILL
XFILL_50_DFFSR_245 gnd vdd FILL
XFILL_12_2_1 gnd vdd FILL
XFILL_65_DFFSR_18 gnd vdd FILL
XFILL_50_DFFSR_256 gnd vdd FILL
XFILL_50_DFFSR_267 gnd vdd FILL
XFILL_65_DFFSR_29 gnd vdd FILL
XFILL_9_AOI21X1_61 gnd vdd FILL
XFILL_9_AOI21X1_72 gnd vdd FILL
XFILL_19_OAI22X1_30 gnd vdd FILL
XFILL_54_DFFSR_200 gnd vdd FILL
XFILL_19_OAI22X1_41 gnd vdd FILL
XFILL_54_DFFSR_211 gnd vdd FILL
XFILL_54_DFFSR_222 gnd vdd FILL
XFILL_54_DFFSR_233 gnd vdd FILL
XFILL_54_DFFSR_244 gnd vdd FILL
XFILL_54_DFFSR_255 gnd vdd FILL
XFILL_3_CLKBUF1_20 gnd vdd FILL
XFILL_54_DFFSR_266 gnd vdd FILL
XFILL_3_CLKBUF1_31 gnd vdd FILL
XFILL_81_DFFSR_100 gnd vdd FILL
XFILL_3_CLKBUF1_42 gnd vdd FILL
XFILL_34_DFFSR_17 gnd vdd FILL
XFILL_81_DFFSR_111 gnd vdd FILL
XFILL_11_MUX2X1_105 gnd vdd FILL
XFILL_58_DFFSR_210 gnd vdd FILL
XFILL_11_MUX2X1_116 gnd vdd FILL
XFILL_81_DFFSR_122 gnd vdd FILL
XFILL_11_MUX2X1_127 gnd vdd FILL
XFILL_34_DFFSR_28 gnd vdd FILL
XFILL_58_DFFSR_221 gnd vdd FILL
XFILL_81_DFFSR_133 gnd vdd FILL
XFILL_34_DFFSR_39 gnd vdd FILL
XFILL_58_DFFSR_232 gnd vdd FILL
XFILL_58_DFFSR_243 gnd vdd FILL
XFILL_81_DFFSR_144 gnd vdd FILL
XFILL_11_MUX2X1_138 gnd vdd FILL
XFILL_11_MUX2X1_149 gnd vdd FILL
XFILL_81_DFFSR_155 gnd vdd FILL
XFILL_58_DFFSR_254 gnd vdd FILL
XFILL_81_DFFSR_166 gnd vdd FILL
XFILL_81_DFFSR_177 gnd vdd FILL
XFILL_58_DFFSR_265 gnd vdd FILL
XFILL_13_CLKBUF1_6 gnd vdd FILL
XFILL_81_DFFSR_188 gnd vdd FILL
XFILL_1_DFFSR_203 gnd vdd FILL
XFILL_12_OAI21X1_10 gnd vdd FILL
XFILL_74_DFFSR_16 gnd vdd FILL
XFILL_85_DFFSR_110 gnd vdd FILL
XFILL_81_DFFSR_199 gnd vdd FILL
XFILL_1_DFFSR_214 gnd vdd FILL
XFILL_74_DFFSR_27 gnd vdd FILL
XFILL_85_DFFSR_121 gnd vdd FILL
XFILL_1_DFFSR_225 gnd vdd FILL
XFILL_12_OAI21X1_21 gnd vdd FILL
XFILL_85_DFFSR_132 gnd vdd FILL
XFILL_1_DFFSR_236 gnd vdd FILL
XFILL_12_OAI21X1_32 gnd vdd FILL
XFILL_74_DFFSR_38 gnd vdd FILL
XFILL_9_5 gnd vdd FILL
XFILL_85_DFFSR_143 gnd vdd FILL
XFILL_1_DFFSR_247 gnd vdd FILL
XFILL_74_DFFSR_49 gnd vdd FILL
XFILL_12_OAI21X1_43 gnd vdd FILL
XFILL_17_MUX2X1_6 gnd vdd FILL
XFILL_85_DFFSR_154 gnd vdd FILL
XFILL_1_DFFSR_258 gnd vdd FILL
XFILL_1_NOR2X1_160 gnd vdd FILL
XFILL_1_DFFSR_269 gnd vdd FILL
XFILL_85_DFFSR_165 gnd vdd FILL
XFILL_1_NOR2X1_171 gnd vdd FILL
XFILL_85_DFFSR_176 gnd vdd FILL
XFILL_17_CLKBUF1_5 gnd vdd FILL
XFILL_5_DFFSR_202 gnd vdd FILL
XFILL_85_DFFSR_187 gnd vdd FILL
XFILL_1_NOR2X1_182 gnd vdd FILL
XFILL_1_NOR2X1_193 gnd vdd FILL
XFILL_2_NAND3X1_2 gnd vdd FILL
XFILL_5_DFFSR_213 gnd vdd FILL
XFILL_85_DFFSR_198 gnd vdd FILL
XFILL_5_DFFSR_224 gnd vdd FILL
XFILL_5_DFFSR_235 gnd vdd FILL
XFILL_8_BUFX4_50 gnd vdd FILL
XFILL_5_DFFSR_246 gnd vdd FILL
XFILL_8_BUFX4_61 gnd vdd FILL
XFILL_43_DFFSR_15 gnd vdd FILL
XFILL_5_DFFSR_257 gnd vdd FILL
XFILL_13_BUFX4_100 gnd vdd FILL
XFILL_5_DFFSR_268 gnd vdd FILL
XFILL_43_DFFSR_26 gnd vdd FILL
XFILL_8_BUFX4_72 gnd vdd FILL
XFILL_8_BUFX4_83 gnd vdd FILL
XFILL_43_DFFSR_37 gnd vdd FILL
XFILL_9_DFFSR_201 gnd vdd FILL
XFILL_8_BUFX4_94 gnd vdd FILL
XFILL_63_6_2 gnd vdd FILL
XFILL_43_DFFSR_48 gnd vdd FILL
XFILL_6_NAND3X1_1 gnd vdd FILL
XFILL_9_DFFSR_212 gnd vdd FILL
XFILL_43_DFFSR_59 gnd vdd FILL
XFILL_9_DFFSR_223 gnd vdd FILL
XFILL_62_1_1 gnd vdd FILL
XFILL_9_DFFSR_234 gnd vdd FILL
XFILL_9_DFFSR_245 gnd vdd FILL
XFILL_9_DFFSR_256 gnd vdd FILL
XFILL_83_DFFSR_14 gnd vdd FILL
XFILL_9_DFFSR_267 gnd vdd FILL
XFILL_83_DFFSR_25 gnd vdd FILL
XFILL_1_MUX2X1_100 gnd vdd FILL
XFILL_83_DFFSR_36 gnd vdd FILL
XFILL_83_DFFSR_47 gnd vdd FILL
XFILL_1_MUX2X1_111 gnd vdd FILL
XFILL_1_MUX2X1_122 gnd vdd FILL
XFILL_83_DFFSR_58 gnd vdd FILL
XFILL_12_DFFSR_14 gnd vdd FILL
XFILL_83_DFFSR_69 gnd vdd FILL
XFILL_12_DFFSR_25 gnd vdd FILL
XFILL_1_MUX2X1_133 gnd vdd FILL
XFILL_1_MUX2X1_144 gnd vdd FILL
XFILL_12_DFFSR_36 gnd vdd FILL
XFILL_1_MUX2X1_155 gnd vdd FILL
XFILL_12_DFFSR_47 gnd vdd FILL
XFILL_87_DFFSR_1 gnd vdd FILL
XFILL_14_NAND3X1_19 gnd vdd FILL
XFILL_12_DFFSR_58 gnd vdd FILL
XFILL_1_MUX2X1_166 gnd vdd FILL
XFILL_12_DFFSR_69 gnd vdd FILL
XFILL_1_MUX2X1_177 gnd vdd FILL
XFILL_1_MUX2X1_188 gnd vdd FILL
XFILL_52_DFFSR_13 gnd vdd FILL
XFILL_34_CLKBUF1_19 gnd vdd FILL
XFILL_21_DFFSR_200 gnd vdd FILL
XFILL_52_DFFSR_24 gnd vdd FILL
XFILL_21_DFFSR_211 gnd vdd FILL
XFILL_52_DFFSR_35 gnd vdd FILL
XFILL_11_NOR2X1_13 gnd vdd FILL
XFILL_21_DFFSR_222 gnd vdd FILL
XFILL_52_DFFSR_46 gnd vdd FILL
XFILL_11_NOR2X1_24 gnd vdd FILL
XFILL_52_DFFSR_57 gnd vdd FILL
XFILL_21_DFFSR_233 gnd vdd FILL
XFILL_11_NOR2X1_35 gnd vdd FILL
XFILL_2_AOI22X1_7 gnd vdd FILL
XFILL_21_DFFSR_244 gnd vdd FILL
XFILL_52_DFFSR_68 gnd vdd FILL
XFILL_11_NOR2X1_46 gnd vdd FILL
XFILL_21_DFFSR_255 gnd vdd FILL
XFILL_52_DFFSR_79 gnd vdd FILL
XFILL_11_NOR2X1_57 gnd vdd FILL
XFILL_11_NOR2X1_68 gnd vdd FILL
XFILL_21_DFFSR_266 gnd vdd FILL
XFILL_11_NOR2X1_79 gnd vdd FILL
XFILL_2_INVX1_206 gnd vdd FILL
XFILL_1_DFFSR_8 gnd vdd FILL
XFILL_9_MUX2X1_5 gnd vdd FILL
XFILL_2_INVX1_217 gnd vdd FILL
XFILL_25_DFFSR_210 gnd vdd FILL
XFILL_2_INVX1_228 gnd vdd FILL
XFILL_25_DFFSR_221 gnd vdd FILL
XFILL_6_AOI22X1_6 gnd vdd FILL
XFILL_21_DFFSR_12 gnd vdd FILL
XFILL_14_DFFSR_6 gnd vdd FILL
XFILL_25_DFFSR_232 gnd vdd FILL
XFILL_25_DFFSR_243 gnd vdd FILL
XFILL_25_DFFSR_254 gnd vdd FILL
XFILL_21_DFFSR_23 gnd vdd FILL
XFILL_71_DFFSR_7 gnd vdd FILL
XFILL_21_DFFSR_34 gnd vdd FILL
XFILL_21_DFFSR_45 gnd vdd FILL
XFILL_25_DFFSR_265 gnd vdd FILL
XFILL_21_DFFSR_56 gnd vdd FILL
XFILL_6_INVX1_205 gnd vdd FILL
XFILL_21_DFFSR_67 gnd vdd FILL
XFILL_6_INVX1_216 gnd vdd FILL
XFILL_52_DFFSR_110 gnd vdd FILL
XFILL_21_DFFSR_78 gnd vdd FILL
XFILL_6_INVX1_227 gnd vdd FILL
XFILL_52_DFFSR_121 gnd vdd FILL
XFILL_21_DFFSR_89 gnd vdd FILL
XFILL_52_DFFSR_132 gnd vdd FILL
XFILL_29_DFFSR_220 gnd vdd FILL
XFILL_61_DFFSR_11 gnd vdd FILL
XFILL_29_DFFSR_231 gnd vdd FILL
XFILL_52_DFFSR_143 gnd vdd FILL
XFILL_29_DFFSR_242 gnd vdd FILL
XFILL_61_DFFSR_22 gnd vdd FILL
XFILL_52_DFFSR_154 gnd vdd FILL
XFILL_29_DFFSR_253 gnd vdd FILL
XFILL_52_DFFSR_165 gnd vdd FILL
XFILL_61_DFFSR_33 gnd vdd FILL
XFILL_29_DFFSR_264 gnd vdd FILL
XFILL_52_DFFSR_176 gnd vdd FILL
XFILL_61_DFFSR_44 gnd vdd FILL
XFILL_29_DFFSR_275 gnd vdd FILL
XFILL_61_DFFSR_55 gnd vdd FILL
XFILL_52_DFFSR_187 gnd vdd FILL
XFILL_61_DFFSR_66 gnd vdd FILL
XFILL_61_DFFSR_77 gnd vdd FILL
XFILL_52_DFFSR_198 gnd vdd FILL
XFILL_56_DFFSR_120 gnd vdd FILL
XFILL_4_NAND3X1_14 gnd vdd FILL
XFILL_56_DFFSR_131 gnd vdd FILL
XFILL_4_NAND3X1_25 gnd vdd FILL
XFILL_61_DFFSR_88 gnd vdd FILL
XFILL_61_DFFSR_99 gnd vdd FILL
XFILL_54_6_2 gnd vdd FILL
XFILL_56_DFFSR_142 gnd vdd FILL
XFILL_4_NAND3X1_36 gnd vdd FILL
XFILL_4_DFFSR_13 gnd vdd FILL
XFILL_56_DFFSR_153 gnd vdd FILL
XFILL_4_NAND3X1_47 gnd vdd FILL
XFILL_4_NAND3X1_58 gnd vdd FILL
XFILL_56_DFFSR_164 gnd vdd FILL
XFILL_4_NAND3X1_69 gnd vdd FILL
XFILL_53_1_1 gnd vdd FILL
XFILL_56_DFFSR_175 gnd vdd FILL
XFILL_4_DFFSR_24 gnd vdd FILL
XFILL_8_NAND2X1_16 gnd vdd FILL
XFILL_4_DFFSR_35 gnd vdd FILL
XFILL_8_NAND2X1_27 gnd vdd FILL
XFILL_56_DFFSR_186 gnd vdd FILL
XFILL_30_DFFSR_10 gnd vdd FILL
XFILL_30_DFFSR_21 gnd vdd FILL
XFILL_4_DFFSR_46 gnd vdd FILL
XFILL_8_NAND2X1_38 gnd vdd FILL
XFILL_8_NAND2X1_49 gnd vdd FILL
XFILL_56_DFFSR_197 gnd vdd FILL
XFILL_4_DFFSR_57 gnd vdd FILL
XFILL_30_DFFSR_32 gnd vdd FILL
XFILL_4_DFFSR_68 gnd vdd FILL
XFILL_30_DFFSR_43 gnd vdd FILL
XFILL_4_DFFSR_79 gnd vdd FILL
XFILL_30_DFFSR_54 gnd vdd FILL
XFILL_30_DFFSR_65 gnd vdd FILL
XFILL_30_DFFSR_76 gnd vdd FILL
XFILL_30_DFFSR_87 gnd vdd FILL
XFILL_30_DFFSR_98 gnd vdd FILL
XFILL_3_DFFSR_101 gnd vdd FILL
XFILL_70_DFFSR_20 gnd vdd FILL
XFILL_3_DFFSR_112 gnd vdd FILL
XFILL_70_DFFSR_31 gnd vdd FILL
XFILL_18_MUX2X1_180 gnd vdd FILL
XFILL_3_DFFSR_123 gnd vdd FILL
XFILL_3_DFFSR_134 gnd vdd FILL
XFILL_70_DFFSR_42 gnd vdd FILL
XFILL_18_MUX2X1_191 gnd vdd FILL
XFILL_3_DFFSR_145 gnd vdd FILL
XFILL_70_DFFSR_53 gnd vdd FILL
XFILL_3_DFFSR_156 gnd vdd FILL
XFILL_70_DFFSR_64 gnd vdd FILL
XFILL_3_DFFSR_167 gnd vdd FILL
XFILL_70_DFFSR_75 gnd vdd FILL
XFILL_3_DFFSR_178 gnd vdd FILL
XFILL_70_DFFSR_86 gnd vdd FILL
XFILL_70_DFFSR_97 gnd vdd FILL
XFILL_7_DFFSR_100 gnd vdd FILL
XFILL_3_DFFSR_189 gnd vdd FILL
XFILL_7_DFFSR_111 gnd vdd FILL
XFILL_38_DFFSR_109 gnd vdd FILL
XFILL_7_DFFSR_122 gnd vdd FILL
XFILL_11_MUX2X1_20 gnd vdd FILL
XFILL_7_DFFSR_133 gnd vdd FILL
XFILL_11_MUX2X1_31 gnd vdd FILL
XFILL_7_DFFSR_144 gnd vdd FILL
XFILL_11_MUX2X1_42 gnd vdd FILL
XFILL_11_MUX2X1_53 gnd vdd FILL
XFILL_7_DFFSR_155 gnd vdd FILL
XDFFSR_180 INVX1_185/A CLKBUF1_34/Y DFFSR_64/R vdd DFFSR_180/D gnd vdd DFFSR
XFILL_11_MUX2X1_64 gnd vdd FILL
XFILL_7_DFFSR_166 gnd vdd FILL
XFILL_7_DFFSR_177 gnd vdd FILL
XFILL_11_MUX2X1_75 gnd vdd FILL
XDFFSR_191 DFFSR_192/D CLKBUF1_7/Y BUFX4_21/Y vdd store gnd vdd DFFSR
XFILL_10_NOR3X1_5 gnd vdd FILL
XFILL_11_MUX2X1_86 gnd vdd FILL
XFILL_7_DFFSR_188 gnd vdd FILL
XFILL_11_MUX2X1_97 gnd vdd FILL
XFILL_7_DFFSR_199 gnd vdd FILL
XFILL_15_MUX2X1_30 gnd vdd FILL
XFILL_15_MUX2X1_41 gnd vdd FILL
XFILL_15_MUX2X1_52 gnd vdd FILL
XFILL_15_MUX2X1_63 gnd vdd FILL
XFILL_3_NOR3X1_12 gnd vdd FILL
XFILL_15_MUX2X1_74 gnd vdd FILL
XFILL_15_MUX2X1_85 gnd vdd FILL
XFILL_3_NOR3X1_23 gnd vdd FILL
XFILL_3_NOR3X1_34 gnd vdd FILL
XFILL_15_MUX2X1_96 gnd vdd FILL
XFILL_3_NOR3X1_45 gnd vdd FILL
XFILL_23_CLKBUF1_15 gnd vdd FILL
XFILL_19_MUX2X1_40 gnd vdd FILL
XFILL_23_CLKBUF1_26 gnd vdd FILL
XFILL_19_MUX2X1_51 gnd vdd FILL
XFILL_23_CLKBUF1_37 gnd vdd FILL
XFILL_19_MUX2X1_62 gnd vdd FILL
XFILL_19_MUX2X1_73 gnd vdd FILL
XFILL_7_NOR3X1_11 gnd vdd FILL
XFILL_19_MUX2X1_84 gnd vdd FILL
XFILL_19_MUX2X1_95 gnd vdd FILL
XFILL_7_NOR3X1_22 gnd vdd FILL
XFILL_6_CLKBUF1_19 gnd vdd FILL
XFILL_0_INVX1_105 gnd vdd FILL
XFILL_7_NOR3X1_33 gnd vdd FILL
XFILL_45_6_2 gnd vdd FILL
XFILL_0_INVX1_116 gnd vdd FILL
XFILL_7_NOR3X1_44 gnd vdd FILL
XFILL_0_INVX1_127 gnd vdd FILL
XFILL_23_DFFSR_120 gnd vdd FILL
XFILL_23_DFFSR_131 gnd vdd FILL
XFILL_1_AOI21X1_16 gnd vdd FILL
XFILL_44_1_1 gnd vdd FILL
XFILL_0_INVX1_138 gnd vdd FILL
XFILL_1_AOI21X1_27 gnd vdd FILL
XFILL_0_INVX1_149 gnd vdd FILL
XFILL_23_DFFSR_142 gnd vdd FILL
XFILL_1_AOI21X1_38 gnd vdd FILL
XFILL_1_AOI21X1_49 gnd vdd FILL
XFILL_23_DFFSR_153 gnd vdd FILL
XFILL_23_DFFSR_164 gnd vdd FILL
XFILL_23_DFFSR_175 gnd vdd FILL
XFILL_11_OAI22X1_18 gnd vdd FILL
XFILL_4_INVX1_104 gnd vdd FILL
XFILL_23_DFFSR_186 gnd vdd FILL
XFILL_11_OAI22X1_29 gnd vdd FILL
XFILL_4_INVX1_115 gnd vdd FILL
XFILL_4_INVX1_126 gnd vdd FILL
XFILL_23_DFFSR_197 gnd vdd FILL
XFILL_4_NOR2X1_104 gnd vdd FILL
XFILL_27_DFFSR_130 gnd vdd FILL
XFILL_4_INVX1_137 gnd vdd FILL
XFILL_4_NOR2X1_115 gnd vdd FILL
XFILL_4_NOR2X1_126 gnd vdd FILL
XFILL_4_INVX1_148 gnd vdd FILL
XFILL_27_DFFSR_141 gnd vdd FILL
XFILL_4_INVX1_159 gnd vdd FILL
XFILL_4_NOR2X1_137 gnd vdd FILL
XFILL_27_DFFSR_152 gnd vdd FILL
XFILL_27_DFFSR_163 gnd vdd FILL
XFILL_4_NOR2X1_148 gnd vdd FILL
XFILL_4_NOR2X1_159 gnd vdd FILL
XFILL_27_DFFSR_174 gnd vdd FILL
XFILL_10_NAND3X1_50 gnd vdd FILL
XFILL_27_DFFSR_185 gnd vdd FILL
XFILL_10_NAND3X1_61 gnd vdd FILL
XFILL_27_DFFSR_196 gnd vdd FILL
XFILL_11_INVX8_4 gnd vdd FILL
XFILL_10_NAND3X1_72 gnd vdd FILL
XFILL_10_NAND3X1_83 gnd vdd FILL
XFILL_2_NOR3X1_4 gnd vdd FILL
XFILL_10_NAND3X1_94 gnd vdd FILL
XFILL_23_NOR3X1_20 gnd vdd FILL
XFILL_23_NOR3X1_31 gnd vdd FILL
XFILL_23_NOR3X1_42 gnd vdd FILL
XFILL_21_MUX2X1_106 gnd vdd FILL
XFILL_21_MUX2X1_117 gnd vdd FILL
XFILL_73_DFFSR_220 gnd vdd FILL
XFILL_21_MUX2X1_128 gnd vdd FILL
XFILL_21_MUX2X1_139 gnd vdd FILL
XFILL_73_DFFSR_231 gnd vdd FILL
XFILL_73_DFFSR_242 gnd vdd FILL
XFILL_73_DFFSR_253 gnd vdd FILL
XFILL_0_DFFSR_50 gnd vdd FILL
XFILL_53_DFFSR_4 gnd vdd FILL
XFILL_73_DFFSR_264 gnd vdd FILL
XFILL_0_DFFSR_61 gnd vdd FILL
XFILL_73_DFFSR_275 gnd vdd FILL
XFILL_0_DFFSR_72 gnd vdd FILL
XFILL_27_NOR3X1_30 gnd vdd FILL
XFILL_0_DFFSR_83 gnd vdd FILL
XFILL_7_2 gnd vdd FILL
XFILL_27_NOR3X1_41 gnd vdd FILL
XFILL_27_NOR3X1_52 gnd vdd FILL
XFILL_9_NOR2X1_204 gnd vdd FILL
XFILL_0_DFFSR_94 gnd vdd FILL
XFILL_77_DFFSR_230 gnd vdd FILL
XFILL_6_OAI22X1_9 gnd vdd FILL
XFILL_1_OAI22X1_13 gnd vdd FILL
XFILL_77_DFFSR_241 gnd vdd FILL
XFILL_1_OAI22X1_24 gnd vdd FILL
XFILL_63_4 gnd vdd FILL
XFILL_1_OAI22X1_35 gnd vdd FILL
XFILL_77_DFFSR_252 gnd vdd FILL
XFILL_1_OAI22X1_46 gnd vdd FILL
XFILL_77_DFFSR_263 gnd vdd FILL
XFILL_32_CLKBUF1_4 gnd vdd FILL
XFILL_77_DFFSR_274 gnd vdd FILL
XFILL_5_OAI21X1_15 gnd vdd FILL
XFILL_56_3 gnd vdd FILL
XFILL_5_OAI21X1_26 gnd vdd FILL
XFILL_5_OAI21X1_37 gnd vdd FILL
XFILL_5_OAI21X1_48 gnd vdd FILL
XFILL_36_6_2 gnd vdd FILL
XFILL_35_1_1 gnd vdd FILL
XFILL_5_DFFSR_9 gnd vdd FILL
XFILL_55_DFFSR_209 gnd vdd FILL
XFILL_18_DFFSR_7 gnd vdd FILL
XFILL_4_NAND2X1_80 gnd vdd FILL
XFILL_75_DFFSR_8 gnd vdd FILL
XFILL_4_NAND2X1_91 gnd vdd FILL
XFILL_9_BUFX4_17 gnd vdd FILL
XFILL_9_BUFX4_28 gnd vdd FILL
XFILL_9_BUFX4_39 gnd vdd FILL
XFILL_12_CLKBUF1_11 gnd vdd FILL
XFILL_12_CLKBUF1_22 gnd vdd FILL
XFILL_82_DFFSR_109 gnd vdd FILL
XFILL_59_DFFSR_208 gnd vdd FILL
XFILL_12_CLKBUF1_33 gnd vdd FILL
XFILL_59_DFFSR_219 gnd vdd FILL
XFILL_86_DFFSR_108 gnd vdd FILL
XFILL_86_DFFSR_119 gnd vdd FILL
XFILL_10_NOR2X1_140 gnd vdd FILL
XFILL_10_NOR2X1_151 gnd vdd FILL
XFILL_10_NOR2X1_162 gnd vdd FILL
XFILL_10_NOR2X1_173 gnd vdd FILL
XFILL_10_NOR2X1_184 gnd vdd FILL
XFILL_40_DFFSR_220 gnd vdd FILL
XFILL_10_NOR2X1_195 gnd vdd FILL
XFILL_40_DFFSR_231 gnd vdd FILL
XFILL_40_DFFSR_242 gnd vdd FILL
XFILL_40_DFFSR_253 gnd vdd FILL
XFILL_40_DFFSR_264 gnd vdd FILL
XNAND3X1_2 INVX2_2/A AND2X2_6/B NAND3X1_2/C gnd OAI22X1_1/B vdd NAND3X1
XFILL_40_DFFSR_275 gnd vdd FILL
XFILL_8_AOI21X1_80 gnd vdd FILL
XFILL_44_DFFSR_230 gnd vdd FILL
XFILL_44_DFFSR_241 gnd vdd FILL
XFILL_44_DFFSR_252 gnd vdd FILL
XFILL_13_BUFX4_11 gnd vdd FILL
XFILL_13_BUFX4_22 gnd vdd FILL
XFILL_44_DFFSR_263 gnd vdd FILL
XFILL_44_DFFSR_274 gnd vdd FILL
XFILL_13_BUFX4_33 gnd vdd FILL
XFILL_27_6_2 gnd vdd FILL
XFILL_12_BUFX4_7 gnd vdd FILL
XFILL_10_MUX2X1_102 gnd vdd FILL
XFILL_2_6_2 gnd vdd FILL
XFILL_13_BUFX4_44 gnd vdd FILL
XFILL_10_MUX2X1_113 gnd vdd FILL
XFILL_13_BUFX4_55 gnd vdd FILL
XFILL_71_DFFSR_130 gnd vdd FILL
XFILL_10_MUX2X1_124 gnd vdd FILL
XFILL_26_1_1 gnd vdd FILL
XFILL_13_BUFX4_66 gnd vdd FILL
XFILL_10_MUX2X1_135 gnd vdd FILL
XFILL_1_1_1 gnd vdd FILL
XFILL_13_BUFX4_77 gnd vdd FILL
XFILL_48_DFFSR_240 gnd vdd FILL
XFILL_13_BUFX4_88 gnd vdd FILL
XFILL_71_DFFSR_141 gnd vdd FILL
XFILL_71_DFFSR_152 gnd vdd FILL
XFILL_10_MUX2X1_146 gnd vdd FILL
XFILL_48_DFFSR_251 gnd vdd FILL
XFILL_13_BUFX4_99 gnd vdd FILL
XFILL_48_DFFSR_262 gnd vdd FILL
XFILL_71_DFFSR_163 gnd vdd FILL
XFILL_10_MUX2X1_157 gnd vdd FILL
XFILL_71_DFFSR_174 gnd vdd FILL
XFILL_10_MUX2X1_168 gnd vdd FILL
XFILL_48_DFFSR_273 gnd vdd FILL
XFILL_71_DFFSR_185 gnd vdd FILL
XFILL_10_MUX2X1_179 gnd vdd FILL
XFILL_71_DFFSR_196 gnd vdd FILL
XFILL_22_DFFSR_209 gnd vdd FILL
XFILL_75_DFFSR_140 gnd vdd FILL
XFILL_11_OAI21X1_40 gnd vdd FILL
XFILL_75_DFFSR_151 gnd vdd FILL
XFILL_75_DFFSR_162 gnd vdd FILL
XFILL_75_DFFSR_173 gnd vdd FILL
XFILL_75_DFFSR_184 gnd vdd FILL
XFILL_75_DFFSR_195 gnd vdd FILL
XFILL_0_NOR2X1_190 gnd vdd FILL
XFILL_10_5_2 gnd vdd FILL
XFILL_26_DFFSR_208 gnd vdd FILL
XAOI22X1_7 NOR2X1_40/Y INVX1_176/A INVX1_171/A NOR2X1_41/Y gnd AOI22X1_7/Y vdd AOI22X1
XFILL_26_DFFSR_219 gnd vdd FILL
XFILL_79_DFFSR_150 gnd vdd FILL
XFILL_7_INVX1_12 gnd vdd FILL
XFILL_79_DFFSR_161 gnd vdd FILL
XFILL_7_INVX1_23 gnd vdd FILL
XFILL_7_INVX1_34 gnd vdd FILL
XINVX1_206 DFFSR_76/Q gnd OAI21X1_5/A vdd INVX1
XFILL_79_DFFSR_172 gnd vdd FILL
XFILL_8_AND2X2_4 gnd vdd FILL
XFILL_79_DFFSR_183 gnd vdd FILL
XFILL_7_INVX1_45 gnd vdd FILL
XINVX1_217 DFFSR_70/Q gnd INVX1_217/Y vdd INVX1
XFILL_7_INVX1_56 gnd vdd FILL
XFILL_79_DFFSR_194 gnd vdd FILL
XFILL_53_DFFSR_108 gnd vdd FILL
XFILL_7_INVX1_67 gnd vdd FILL
XINVX1_228 DFFSR_54/Q gnd OAI22X1_5/A vdd INVX1
XFILL_53_DFFSR_119 gnd vdd FILL
XFILL_7_INVX1_78 gnd vdd FILL
XFILL_7_INVX1_89 gnd vdd FILL
XFILL_9_2_1 gnd vdd FILL
XFILL_57_DFFSR_107 gnd vdd FILL
XFILL_57_DFFSR_118 gnd vdd FILL
XFILL_0_MUX2X1_130 gnd vdd FILL
XFILL_0_MUX2X1_141 gnd vdd FILL
XFILL_57_DFFSR_129 gnd vdd FILL
XFILL_35_DFFSR_1 gnd vdd FILL
XFILL_5_BUFX4_10 gnd vdd FILL
XFILL_0_MUX2X1_152 gnd vdd FILL
XFILL_0_MUX2X1_163 gnd vdd FILL
XFILL_5_BUFX4_21 gnd vdd FILL
XFILL_13_NAND3X1_16 gnd vdd FILL
XFILL_5_BUFX4_32 gnd vdd FILL
XNAND2X1_17 NAND3X1_67/Y OAI21X1_23/Y gnd NOR3X1_9/B vdd NAND2X1
XFILL_5_BUFX4_43 gnd vdd FILL
XNAND2X1_28 BUFX4_89/Y NOR2X1_44/Y gnd NOR2X1_98/B vdd NAND2X1
XFILL_13_NAND3X1_27 gnd vdd FILL
XFILL_0_MUX2X1_174 gnd vdd FILL
XFILL_0_MUX2X1_185 gnd vdd FILL
XFILL_5_BUFX4_54 gnd vdd FILL
XFILL_13_NAND3X1_38 gnd vdd FILL
XNAND2X1_39 AND2X2_1/B AND2X2_6/A gnd NOR3X1_29/B vdd NAND2X1
XFILL_13_NAND3X1_49 gnd vdd FILL
XFILL_40_DFFSR_19 gnd vdd FILL
XFILL_5_BUFX4_65 gnd vdd FILL
XFILL_5_BUFX4_76 gnd vdd FILL
XFILL_33_CLKBUF1_16 gnd vdd FILL
XFILL_5_BUFX4_87 gnd vdd FILL
XFILL_33_CLKBUF1_27 gnd vdd FILL
XFILL_5_BUFX4_98 gnd vdd FILL
XFILL_33_CLKBUF1_38 gnd vdd FILL
XFILL_11_DFFSR_230 gnd vdd FILL
XFILL_11_DFFSR_241 gnd vdd FILL
XFILL_18_6_2 gnd vdd FILL
XFILL_11_DFFSR_252 gnd vdd FILL
XFILL_17_1_1 gnd vdd FILL
XFILL_11_DFFSR_263 gnd vdd FILL
XFILL_11_DFFSR_274 gnd vdd FILL
XFILL_80_DFFSR_18 gnd vdd FILL
XFILL_80_DFFSR_29 gnd vdd FILL
XFILL_23_MUX2X1_8 gnd vdd FILL
XFILL_15_DFFSR_240 gnd vdd FILL
XFILL_60_4_2 gnd vdd FILL
XFILL_15_DFFSR_251 gnd vdd FILL
XFILL_28_7 gnd vdd FILL
XFILL_57_DFFSR_5 gnd vdd FILL
XFILL_15_DFFSR_262 gnd vdd FILL
XFILL_8_DFFSR_109 gnd vdd FILL
XFILL_15_DFFSR_273 gnd vdd FILL
XFILL_12_MUX2X1_18 gnd vdd FILL
XFILL_12_MUX2X1_29 gnd vdd FILL
XFILL_42_DFFSR_140 gnd vdd FILL
XFILL_3_AOI21X1_5 gnd vdd FILL
XFILL_42_DFFSR_151 gnd vdd FILL
XFILL_19_DFFSR_250 gnd vdd FILL
XFILL_42_DFFSR_162 gnd vdd FILL
XFILL_19_DFFSR_261 gnd vdd FILL
XFILL_42_DFFSR_173 gnd vdd FILL
XFILL_42_DFFSR_184 gnd vdd FILL
XFILL_19_DFFSR_272 gnd vdd FILL
XFILL_16_MUX2X1_17 gnd vdd FILL
XFILL_42_DFFSR_195 gnd vdd FILL
XFILL_16_MUX2X1_28 gnd vdd FILL
XFILL_3_NAND3X1_11 gnd vdd FILL
XFILL_16_MUX2X1_39 gnd vdd FILL
XFILL_3_NAND3X1_22 gnd vdd FILL
XFILL_7_AOI21X1_4 gnd vdd FILL
XFILL_3_NAND3X1_33 gnd vdd FILL
XFILL_6_MUX2X1_9 gnd vdd FILL
XFILL_46_DFFSR_150 gnd vdd FILL
XFILL_3_NAND3X1_44 gnd vdd FILL
XNOR3X1_5 NOR3X1_5/A NOR3X1_5/B NOR3X1_5/C gnd NOR3X1_7/A vdd NOR3X1
XFILL_46_DFFSR_161 gnd vdd FILL
XFILL_3_NAND3X1_55 gnd vdd FILL
XFILL_3_NAND3X1_66 gnd vdd FILL
XFILL_46_DFFSR_172 gnd vdd FILL
XFILL_7_NAND2X1_13 gnd vdd FILL
XFILL_3_NAND3X1_77 gnd vdd FILL
XFILL_46_DFFSR_183 gnd vdd FILL
XFILL_7_NAND2X1_24 gnd vdd FILL
XFILL_46_DFFSR_194 gnd vdd FILL
XFILL_7_NAND2X1_35 gnd vdd FILL
XFILL_20_DFFSR_108 gnd vdd FILL
XFILL_3_NAND3X1_88 gnd vdd FILL
XFILL_7_NAND2X1_46 gnd vdd FILL
XFILL_3_NAND3X1_99 gnd vdd FILL
XFILL_7_NAND2X1_57 gnd vdd FILL
XFILL_20_DFFSR_119 gnd vdd FILL
XFILL_7_NAND2X1_68 gnd vdd FILL
XFILL_79_DFFSR_9 gnd vdd FILL
XFILL_7_NAND2X1_79 gnd vdd FILL
XFILL_12_AOI22X1_1 gnd vdd FILL
XFILL_24_DFFSR_107 gnd vdd FILL
XFILL_24_DFFSR_118 gnd vdd FILL
XFILL_24_DFFSR_129 gnd vdd FILL
XFILL_61_1 gnd vdd FILL
XFILL_10_AOI21X1_18 gnd vdd FILL
XFILL_10_AOI21X1_29 gnd vdd FILL
XFILL_1_DFFSR_17 gnd vdd FILL
XFILL_28_DFFSR_106 gnd vdd FILL
XFILL_28_DFFSR_117 gnd vdd FILL
XFILL_1_DFFSR_28 gnd vdd FILL
XFILL_11_NOR2X1_5 gnd vdd FILL
XFILL_1_DFFSR_39 gnd vdd FILL
XFILL_28_DFFSR_128 gnd vdd FILL
XFILL_28_DFFSR_139 gnd vdd FILL
XFILL_3_INVX1_60 gnd vdd FILL
XFILL_7_AOI22X1_11 gnd vdd FILL
XFILL_3_INVX1_71 gnd vdd FILL
XFILL_20_NOR3X1_19 gnd vdd FILL
XFILL_3_INVX1_82 gnd vdd FILL
XFILL_51_4_2 gnd vdd FILL
XFILL_3_INVX1_93 gnd vdd FILL
XFILL_49_DFFSR_30 gnd vdd FILL
XFILL_70_DFFSR_208 gnd vdd FILL
XFILL_49_DFFSR_41 gnd vdd FILL
XFILL_70_DFFSR_219 gnd vdd FILL
XFILL_49_DFFSR_52 gnd vdd FILL
XFILL_49_DFFSR_63 gnd vdd FILL
XFILL_10_MUX2X1_3 gnd vdd FILL
XFILL_49_DFFSR_74 gnd vdd FILL
XFILL_49_DFFSR_85 gnd vdd FILL
XFILL_24_NOR3X1_18 gnd vdd FILL
XFILL_49_DFFSR_96 gnd vdd FILL
XFILL_24_NOR3X1_29 gnd vdd FILL
XFILL_22_CLKBUF1_12 gnd vdd FILL
XFILL_74_DFFSR_207 gnd vdd FILL
XFILL_22_CLKBUF1_23 gnd vdd FILL
XFILL_22_CLKBUF1_34 gnd vdd FILL
XFILL_74_DFFSR_218 gnd vdd FILL
XFILL_74_DFFSR_229 gnd vdd FILL
XFILL_18_DFFSR_40 gnd vdd FILL
XFILL_28_NOR3X1_17 gnd vdd FILL
XFILL_1_BUFX4_80 gnd vdd FILL
XFILL_18_DFFSR_51 gnd vdd FILL
XFILL_5_CLKBUF1_16 gnd vdd FILL
XFILL_1_BUFX4_91 gnd vdd FILL
XFILL_28_NOR3X1_28 gnd vdd FILL
XFILL_18_DFFSR_62 gnd vdd FILL
XFILL_5_CLKBUF1_27 gnd vdd FILL
XFILL_5_CLKBUF1_38 gnd vdd FILL
XFILL_28_NOR3X1_39 gnd vdd FILL
XFILL_78_DFFSR_206 gnd vdd FILL
XFILL_18_DFFSR_73 gnd vdd FILL
XFILL_18_DFFSR_84 gnd vdd FILL
XFILL_0_AOI21X1_13 gnd vdd FILL
XFILL_18_DFFSR_95 gnd vdd FILL
XFILL_78_DFFSR_217 gnd vdd FILL
XFILL_0_AOI21X1_24 gnd vdd FILL
XFILL_78_DFFSR_228 gnd vdd FILL
XFILL_0_AOI21X1_35 gnd vdd FILL
XFILL_0_AOI21X1_46 gnd vdd FILL
XFILL_13_DFFSR_150 gnd vdd FILL
XFILL_78_DFFSR_239 gnd vdd FILL
XFILL_13_DFFSR_161 gnd vdd FILL
XFILL_0_AOI21X1_57 gnd vdd FILL
XFILL_29_NOR3X1_3 gnd vdd FILL
XFILL_13_DFFSR_172 gnd vdd FILL
XFILL_2_CLKBUF1_4 gnd vdd FILL
XFILL_10_OAI22X1_15 gnd vdd FILL
XFILL_0_AOI21X1_68 gnd vdd FILL
XFILL_13_DFFSR_183 gnd vdd FILL
XFILL_10_OAI22X1_26 gnd vdd FILL
XFILL_58_DFFSR_50 gnd vdd FILL
XFILL_13_DFFSR_194 gnd vdd FILL
XFILL_0_AOI21X1_79 gnd vdd FILL
XFILL_10_OAI22X1_37 gnd vdd FILL
XFILL_58_DFFSR_61 gnd vdd FILL
XFILL_58_DFFSR_72 gnd vdd FILL
XFILL_3_NOR2X1_101 gnd vdd FILL
XFILL_10_OAI22X1_48 gnd vdd FILL
XFILL_58_DFFSR_83 gnd vdd FILL
XFILL_14_OAI21X1_17 gnd vdd FILL
XFILL_3_NOR2X1_112 gnd vdd FILL
XFILL_3_NOR2X1_123 gnd vdd FILL
XFILL_58_DFFSR_94 gnd vdd FILL
XFILL_3_NOR2X1_134 gnd vdd FILL
XFILL_14_OAI21X1_28 gnd vdd FILL
XFILL_3_NOR2X1_145 gnd vdd FILL
XFILL_14_OAI21X1_39 gnd vdd FILL
XFILL_17_DFFSR_160 gnd vdd FILL
XFILL_59_5_2 gnd vdd FILL
XFILL_6_CLKBUF1_3 gnd vdd FILL
XFILL_3_NOR2X1_156 gnd vdd FILL
XFILL_17_DFFSR_171 gnd vdd FILL
XFILL_3_NOR2X1_4 gnd vdd FILL
XFILL_3_NOR2X1_167 gnd vdd FILL
XFILL_17_DFFSR_182 gnd vdd FILL
XFILL_58_0_1 gnd vdd FILL
XFILL_3_NOR2X1_178 gnd vdd FILL
XFILL_17_DFFSR_193 gnd vdd FILL
XFILL_3_NOR2X1_189 gnd vdd FILL
XFILL_27_DFFSR_60 gnd vdd FILL
XFILL_27_DFFSR_71 gnd vdd FILL
XFILL_27_DFFSR_82 gnd vdd FILL
XFILL_27_DFFSR_93 gnd vdd FILL
XFILL_13_NOR3X1_50 gnd vdd FILL
XFILL_20_MUX2X1_103 gnd vdd FILL
XFILL_2_MUX2X1_2 gnd vdd FILL
XFILL_20_MUX2X1_114 gnd vdd FILL
XFILL_20_MUX2X1_125 gnd vdd FILL
XFILL_67_DFFSR_70 gnd vdd FILL
XFILL_20_MUX2X1_136 gnd vdd FILL
XFILL_42_4_2 gnd vdd FILL
XFILL_67_DFFSR_81 gnd vdd FILL
XFILL_67_DFFSR_92 gnd vdd FILL
XFILL_63_DFFSR_250 gnd vdd FILL
XFILL_20_MUX2X1_147 gnd vdd FILL
XFILL_20_MUX2X1_158 gnd vdd FILL
XFILL_63_DFFSR_261 gnd vdd FILL
XFILL_20_MUX2X1_169 gnd vdd FILL
XFILL_3_MUX2X1_107 gnd vdd FILL
XFILL_63_DFFSR_272 gnd vdd FILL
XFILL_3_MUX2X1_118 gnd vdd FILL
XFILL_3_MUX2X1_129 gnd vdd FILL
XFILL_39_DFFSR_2 gnd vdd FILL
XFILL_8_NOR2X1_201 gnd vdd FILL
XFILL_0_OAI22X1_10 gnd vdd FILL
XFILL_0_OAI22X1_21 gnd vdd FILL
XFILL_0_OAI22X1_32 gnd vdd FILL
XFILL_0_OAI22X1_43 gnd vdd FILL
XFILL_67_DFFSR_260 gnd vdd FILL
XFILL_67_DFFSR_271 gnd vdd FILL
XFILL_22_CLKBUF1_1 gnd vdd FILL
XFILL_4_OAI21X1_12 gnd vdd FILL
XFILL_36_DFFSR_80 gnd vdd FILL
XFILL_4_OAI21X1_23 gnd vdd FILL
XFILL_36_DFFSR_91 gnd vdd FILL
XFILL_0_NOR2X1_11 gnd vdd FILL
XFILL_4_OAI21X1_34 gnd vdd FILL
XFILL_41_DFFSR_207 gnd vdd FILL
XFILL_0_NOR2X1_22 gnd vdd FILL
XFILL_0_NOR2X1_33 gnd vdd FILL
XFILL_41_DFFSR_218 gnd vdd FILL
XFILL_4_OAI21X1_45 gnd vdd FILL
XFILL_0_NOR2X1_44 gnd vdd FILL
XFILL_3_OAI21X1_8 gnd vdd FILL
XFILL_41_DFFSR_229 gnd vdd FILL
XFILL_0_NOR2X1_55 gnd vdd FILL
XAOI21X1_70 INVX1_82/A INVX1_127/Y OAI22X1_6/Y gnd NAND3X1_84/A vdd AOI21X1
XFILL_0_NOR2X1_66 gnd vdd FILL
XAOI21X1_81 BUFX4_68/Y AOI21X1_3/B NOR2X1_125/Y gnd DFFSR_149/D vdd AOI21X1
XFILL_0_NOR2X1_77 gnd vdd FILL
XFILL_0_NOR2X1_88 gnd vdd FILL
XFILL_45_DFFSR_206 gnd vdd FILL
XFILL_76_DFFSR_90 gnd vdd FILL
XFILL_0_NOR2X1_99 gnd vdd FILL
XFILL_4_NOR2X1_10 gnd vdd FILL
XFILL_23_DFFSR_8 gnd vdd FILL
XFILL_4_NOR2X1_21 gnd vdd FILL
XFILL_45_DFFSR_217 gnd vdd FILL
XFILL_7_OAI21X1_7 gnd vdd FILL
XFILL_4_NOR2X1_32 gnd vdd FILL
XFILL_80_DFFSR_9 gnd vdd FILL
XFILL_4_NOR2X1_43 gnd vdd FILL
XFILL_45_DFFSR_228 gnd vdd FILL
XFILL_45_DFFSR_239 gnd vdd FILL
XFILL_4_NOR2X1_54 gnd vdd FILL
XFILL_4_NOR2X1_65 gnd vdd FILL
XFILL_4_NOR2X1_76 gnd vdd FILL
XFILL_4_NOR2X1_87 gnd vdd FILL
XFILL_4_NOR2X1_98 gnd vdd FILL
XFILL_72_DFFSR_106 gnd vdd FILL
XFILL_49_DFFSR_205 gnd vdd FILL
XFILL_11_CLKBUF1_30 gnd vdd FILL
XFILL_49_DFFSR_216 gnd vdd FILL
XFILL_72_DFFSR_117 gnd vdd FILL
XFILL_8_NOR2X1_20 gnd vdd FILL
XFILL_11_CLKBUF1_41 gnd vdd FILL
XFILL_8_NOR2X1_31 gnd vdd FILL
XFILL_72_DFFSR_128 gnd vdd FILL
XFILL_49_0_1 gnd vdd FILL
XFILL_8_NOR2X1_42 gnd vdd FILL
XFILL_49_DFFSR_227 gnd vdd FILL
XFILL_72_DFFSR_139 gnd vdd FILL
XFILL_8_NOR2X1_53 gnd vdd FILL
XFILL_12_OAI22X1_4 gnd vdd FILL
XFILL_49_DFFSR_238 gnd vdd FILL
XFILL_49_DFFSR_249 gnd vdd FILL
XFILL_8_NOR2X1_64 gnd vdd FILL
XFILL_8_NOR2X1_75 gnd vdd FILL
XFILL_8_NOR2X1_86 gnd vdd FILL
XFILL_8_NOR2X1_97 gnd vdd FILL
XFILL_76_DFFSR_105 gnd vdd FILL
XFILL_76_DFFSR_116 gnd vdd FILL
XFILL_76_DFFSR_127 gnd vdd FILL
XFILL_76_DFFSR_138 gnd vdd FILL
XFILL_16_OAI22X1_3 gnd vdd FILL
XFILL_76_DFFSR_149 gnd vdd FILL
XFILL_61_7_0 gnd vdd FILL
XFILL_33_4_2 gnd vdd FILL
XFILL_26_4 gnd vdd FILL
XFILL_30_DFFSR_250 gnd vdd FILL
XFILL_19_3 gnd vdd FILL
XFILL_30_DFFSR_261 gnd vdd FILL
XFILL_30_DFFSR_272 gnd vdd FILL
XFILL_34_DFFSR_260 gnd vdd FILL
XFILL_34_DFFSR_271 gnd vdd FILL
XFILL_4_NAND2X1_9 gnd vdd FILL
XFILL_0_MUX2X1_40 gnd vdd FILL
XFILL_0_MUX2X1_51 gnd vdd FILL
XFILL_0_MUX2X1_62 gnd vdd FILL
XFILL_0_MUX2X1_73 gnd vdd FILL
XFILL_0_MUX2X1_84 gnd vdd FILL
XFILL_61_DFFSR_160 gnd vdd FILL
XFILL_0_MUX2X1_95 gnd vdd FILL
XFILL_38_DFFSR_270 gnd vdd FILL
XFILL_61_DFFSR_171 gnd vdd FILL
XFILL_61_DFFSR_182 gnd vdd FILL
XFILL_61_DFFSR_193 gnd vdd FILL
XFILL_8_NAND2X1_8 gnd vdd FILL
XFILL_12_DFFSR_206 gnd vdd FILL
XFILL_4_MUX2X1_50 gnd vdd FILL
XFILL_12_DFFSR_217 gnd vdd FILL
XFILL_12_DFFSR_228 gnd vdd FILL
XFILL_4_MUX2X1_61 gnd vdd FILL
XFILL_12_DFFSR_239 gnd vdd FILL
XFILL_4_MUX2X1_72 gnd vdd FILL
XFILL_4_MUX2X1_83 gnd vdd FILL
XFILL_4_MUX2X1_94 gnd vdd FILL
XFILL_65_DFFSR_170 gnd vdd FILL
XFILL_65_DFFSR_181 gnd vdd FILL
XFILL_65_DFFSR_192 gnd vdd FILL
XFILL_16_DFFSR_205 gnd vdd FILL
XFILL_10_BUFX4_15 gnd vdd FILL
XFILL_13_NAND3X1_5 gnd vdd FILL
XFILL_10_BUFX4_26 gnd vdd FILL
XFILL_16_DFFSR_216 gnd vdd FILL
XFILL_10_BUFX4_37 gnd vdd FILL
XFILL_8_MUX2X1_60 gnd vdd FILL
XFILL_16_DFFSR_227 gnd vdd FILL
XFILL_8_MUX2X1_71 gnd vdd FILL
XFILL_10_BUFX4_48 gnd vdd FILL
XFILL_16_DFFSR_238 gnd vdd FILL
XFILL_10_BUFX4_59 gnd vdd FILL
XFILL_16_DFFSR_249 gnd vdd FILL
XFILL_8_MUX2X1_82 gnd vdd FILL
XFILL_8_MUX2X1_93 gnd vdd FILL
XFILL_69_DFFSR_180 gnd vdd FILL
XFILL_69_DFFSR_191 gnd vdd FILL
XFILL_43_DFFSR_105 gnd vdd FILL
XFILL_43_DFFSR_116 gnd vdd FILL
XFILL_43_DFFSR_127 gnd vdd FILL
XFILL_43_DFFSR_138 gnd vdd FILL
XFILL_43_DFFSR_149 gnd vdd FILL
XFILL_52_7_0 gnd vdd FILL
XFILL_24_4_2 gnd vdd FILL
XFILL_47_DFFSR_104 gnd vdd FILL
XFILL_47_DFFSR_115 gnd vdd FILL
XFILL_40_DFFSR_2 gnd vdd FILL
XFILL_47_DFFSR_126 gnd vdd FILL
XFILL_8_DFFSR_1 gnd vdd FILL
XFILL_47_DFFSR_137 gnd vdd FILL
XFILL_47_DFFSR_148 gnd vdd FILL
XFILL_12_NAND3X1_13 gnd vdd FILL
XFILL_20_MUX2X1_70 gnd vdd FILL
XFILL_47_DFFSR_159 gnd vdd FILL
XFILL_12_NAND3X1_24 gnd vdd FILL
XFILL_20_MUX2X1_81 gnd vdd FILL
XFILL_12_NAND3X1_35 gnd vdd FILL
XFILL_20_MUX2X1_92 gnd vdd FILL
XFILL_4_INVX1_16 gnd vdd FILL
XFILL_12_NAND3X1_46 gnd vdd FILL
XFILL_12_NAND3X1_57 gnd vdd FILL
XFILL_12_NAND3X1_68 gnd vdd FILL
XFILL_4_INVX1_27 gnd vdd FILL
XFILL_4_INVX1_38 gnd vdd FILL
XFILL_32_CLKBUF1_13 gnd vdd FILL
XFILL_32_CLKBUF1_24 gnd vdd FILL
XFILL_12_NAND3X1_79 gnd vdd FILL
XFILL_5_AND2X2_8 gnd vdd FILL
XFILL_4_INVX1_49 gnd vdd FILL
XFILL_32_CLKBUF1_35 gnd vdd FILL
XFILL_3_BUFX2_7 gnd vdd FILL
XFILL_17_AOI22X1_9 gnd vdd FILL
XFILL_2_BUFX4_14 gnd vdd FILL
XFILL_62_DFFSR_6 gnd vdd FILL
XFILL_2_BUFX4_25 gnd vdd FILL
XFILL_2_BUFX4_36 gnd vdd FILL
XFILL_2_BUFX4_47 gnd vdd FILL
XFILL_19_DFFSR_18 gnd vdd FILL
XFILL_2_BUFX4_58 gnd vdd FILL
XFILL_7_5_2 gnd vdd FILL
XFILL_19_DFFSR_29 gnd vdd FILL
XFILL_2_BUFX4_69 gnd vdd FILL
XFILL_14_OR2X2_1 gnd vdd FILL
XFILL_6_0_1 gnd vdd FILL
XFILL_32_DFFSR_170 gnd vdd FILL
XFILL_32_DFFSR_181 gnd vdd FILL
XFILL_32_DFFSR_192 gnd vdd FILL
XFILL_59_DFFSR_17 gnd vdd FILL
XFILL_59_DFFSR_28 gnd vdd FILL
XFILL_59_DFFSR_39 gnd vdd FILL
XFILL_2_NAND3X1_30 gnd vdd FILL
XFILL_2_NAND3X1_41 gnd vdd FILL
XFILL_6_NAND2X1_10 gnd vdd FILL
XFILL_2_NAND3X1_52 gnd vdd FILL
XFILL_2_NAND3X1_63 gnd vdd FILL
XFILL_36_DFFSR_180 gnd vdd FILL
XFILL_2_NAND3X1_74 gnd vdd FILL
XFILL_6_NAND2X1_21 gnd vdd FILL
XFILL_2_NAND3X1_85 gnd vdd FILL
XFILL_6_NAND2X1_32 gnd vdd FILL
XFILL_36_DFFSR_191 gnd vdd FILL
XFILL_10_DFFSR_105 gnd vdd FILL
XFILL_43_7_0 gnd vdd FILL
XFILL_2_BUFX4_1 gnd vdd FILL
XFILL_6_NAND2X1_43 gnd vdd FILL
XFILL_2_NAND3X1_96 gnd vdd FILL
XFILL_10_DFFSR_116 gnd vdd FILL
XFILL_15_4_2 gnd vdd FILL
XFILL_6_NAND2X1_54 gnd vdd FILL
XFILL_27_DFFSR_9 gnd vdd FILL
XFILL_6_NAND2X1_65 gnd vdd FILL
XFILL_10_DFFSR_127 gnd vdd FILL
XFILL_10_DFFSR_138 gnd vdd FILL
XFILL_28_DFFSR_16 gnd vdd FILL
XFILL_6_NAND2X1_76 gnd vdd FILL
XFILL_10_DFFSR_149 gnd vdd FILL
XFILL_6_NAND2X1_87 gnd vdd FILL
XMUX2X1_3 MUX2X1_7/B MUX2X1_3/B MUX2X1_3/S gnd MUX2X1_3/Y vdd MUX2X1
XFILL_28_DFFSR_27 gnd vdd FILL
XFILL_28_DFFSR_38 gnd vdd FILL
XFILL_28_DFFSR_49 gnd vdd FILL
XFILL_14_DFFSR_104 gnd vdd FILL
XFILL_14_CLKBUF1_18 gnd vdd FILL
XFILL_14_DFFSR_115 gnd vdd FILL
XFILL_14_CLKBUF1_29 gnd vdd FILL
XFILL_14_DFFSR_126 gnd vdd FILL
XFILL_14_DFFSR_137 gnd vdd FILL
XFILL_68_DFFSR_15 gnd vdd FILL
XFILL_14_DFFSR_148 gnd vdd FILL
XFILL_68_DFFSR_26 gnd vdd FILL
XFILL_14_DFFSR_159 gnd vdd FILL
XFILL_68_DFFSR_37 gnd vdd FILL
XFILL_68_DFFSR_48 gnd vdd FILL
XFILL_68_DFFSR_59 gnd vdd FILL
XFILL_82_DFFSR_270 gnd vdd FILL
XFILL_18_DFFSR_103 gnd vdd FILL
XFILL_18_DFFSR_114 gnd vdd FILL
XFILL_1_INVX1_5 gnd vdd FILL
XFILL_18_DFFSR_125 gnd vdd FILL
XFILL_18_DFFSR_136 gnd vdd FILL
XFILL_18_DFFSR_147 gnd vdd FILL
XFILL_18_DFFSR_158 gnd vdd FILL
XCLKBUF1_4 BUFX4_9/Y gnd CLKBUF1_4/Y vdd CLKBUF1
XFILL_18_DFFSR_169 gnd vdd FILL
XFILL_10_NOR3X1_16 gnd vdd FILL
XFILL_37_DFFSR_14 gnd vdd FILL
XFILL_10_NOR3X1_27 gnd vdd FILL
XFILL_37_DFFSR_25 gnd vdd FILL
XFILL_37_DFFSR_36 gnd vdd FILL
XFILL_10_NOR3X1_38 gnd vdd FILL
XFILL_10_NOR3X1_49 gnd vdd FILL
XFILL_60_DFFSR_205 gnd vdd FILL
XFILL_37_DFFSR_47 gnd vdd FILL
XFILL_37_DFFSR_58 gnd vdd FILL
XFILL_60_DFFSR_216 gnd vdd FILL
XFILL_60_DFFSR_227 gnd vdd FILL
XFILL_37_DFFSR_69 gnd vdd FILL
XFILL_60_DFFSR_238 gnd vdd FILL
XFILL_60_DFFSR_249 gnd vdd FILL
XFILL_14_NOR3X1_15 gnd vdd FILL
XFILL_77_DFFSR_13 gnd vdd FILL
XFILL_14_NOR3X1_26 gnd vdd FILL
XFILL_77_DFFSR_24 gnd vdd FILL
XFILL_77_DFFSR_35 gnd vdd FILL
XFILL_14_NOR3X1_37 gnd vdd FILL
XFILL_21_CLKBUF1_20 gnd vdd FILL
XFILL_77_DFFSR_46 gnd vdd FILL
XFILL_14_NOR3X1_48 gnd vdd FILL
XFILL_64_DFFSR_204 gnd vdd FILL
XFILL_64_DFFSR_215 gnd vdd FILL
XFILL_21_CLKBUF1_31 gnd vdd FILL
XFILL_2_INVX4_1 gnd vdd FILL
XFILL_77_DFFSR_57 gnd vdd FILL
XFILL_21_CLKBUF1_42 gnd vdd FILL
XFILL_77_DFFSR_68 gnd vdd FILL
XFILL_64_DFFSR_226 gnd vdd FILL
XFILL_64_DFFSR_237 gnd vdd FILL
XFILL_77_DFFSR_79 gnd vdd FILL
XFILL_65_3_2 gnd vdd FILL
XFILL_64_DFFSR_248 gnd vdd FILL
XFILL_0_INVX1_20 gnd vdd FILL
XFILL_18_NOR3X1_14 gnd vdd FILL
XFILL_0_INVX1_31 gnd vdd FILL
XFILL_4_CLKBUF1_13 gnd vdd FILL
XFILL_64_DFFSR_259 gnd vdd FILL
XFILL_18_NOR3X1_25 gnd vdd FILL
XFILL_4_CLKBUF1_24 gnd vdd FILL
XFILL_0_INVX1_42 gnd vdd FILL
XFILL_1_AND2X2_1 gnd vdd FILL
XNOR2X1_202 DFFSR_9/Q NOR2X1_202/B gnd NOR2X1_202/Y vdd NOR2X1
XFILL_18_NOR3X1_36 gnd vdd FILL
XFILL_0_INVX1_53 gnd vdd FILL
XFILL_4_CLKBUF1_35 gnd vdd FILL
XFILL_18_NOR3X1_47 gnd vdd FILL
XFILL_0_INVX1_64 gnd vdd FILL
XFILL_68_DFFSR_203 gnd vdd FILL
XFILL_12_MUX2X1_109 gnd vdd FILL
XFILL_0_INVX1_75 gnd vdd FILL
XFILL_68_DFFSR_214 gnd vdd FILL
XFILL_0_INVX1_86 gnd vdd FILL
XFILL_46_DFFSR_12 gnd vdd FILL
XFILL_46_DFFSR_23 gnd vdd FILL
XFILL_68_DFFSR_225 gnd vdd FILL
XFILL_0_INVX1_97 gnd vdd FILL
XFILL_34_7_0 gnd vdd FILL
XFILL_68_DFFSR_236 gnd vdd FILL
XFILL_46_DFFSR_34 gnd vdd FILL
XFILL_31_2 gnd vdd FILL
XFILL_17_NOR3X1_9 gnd vdd FILL
XFILL_68_DFFSR_247 gnd vdd FILL
XFILL_46_DFFSR_45 gnd vdd FILL
XFILL_46_DFFSR_56 gnd vdd FILL
XFILL_68_DFFSR_258 gnd vdd FILL
XFILL_68_DFFSR_269 gnd vdd FILL
XFILL_46_DFFSR_67 gnd vdd FILL
XFILL_46_DFFSR_78 gnd vdd FILL
XFILL_24_1 gnd vdd FILL
XFILL_46_DFFSR_89 gnd vdd FILL
XFILL_13_OAI21X1_14 gnd vdd FILL
XFILL_86_DFFSR_11 gnd vdd FILL
XFILL_13_OAI21X1_25 gnd vdd FILL
XFILL_2_NOR2X1_120 gnd vdd FILL
XFILL_86_DFFSR_22 gnd vdd FILL
XFILL_2_NOR2X1_131 gnd vdd FILL
XFILL_13_OAI21X1_36 gnd vdd FILL
XFILL_86_DFFSR_33 gnd vdd FILL
XFILL_2_NOR2X1_142 gnd vdd FILL
XFILL_2_NOR2X1_153 gnd vdd FILL
XFILL_13_OAI21X1_47 gnd vdd FILL
XFILL_86_DFFSR_44 gnd vdd FILL
XFILL_86_DFFSR_55 gnd vdd FILL
XFILL_15_DFFSR_11 gnd vdd FILL
XFILL_86_DFFSR_66 gnd vdd FILL
XFILL_2_NOR2X1_164 gnd vdd FILL
XFILL_27_CLKBUF1_9 gnd vdd FILL
XFILL_2_NOR2X1_175 gnd vdd FILL
XFILL_15_DFFSR_22 gnd vdd FILL
XFILL_86_DFFSR_77 gnd vdd FILL
XFILL_15_DFFSR_33 gnd vdd FILL
XFILL_2_NOR2X1_186 gnd vdd FILL
XFILL_2_NOR2X1_197 gnd vdd FILL
XFILL_86_DFFSR_88 gnd vdd FILL
XFILL_15_DFFSR_44 gnd vdd FILL
XFILL_5_NOR2X1_19 gnd vdd FILL
XFILL_15_DFFSR_55 gnd vdd FILL
XFILL_86_DFFSR_99 gnd vdd FILL
XFILL_15_DFFSR_66 gnd vdd FILL
XFILL_26_11 gnd vdd FILL
XFILL_15_DFFSR_77 gnd vdd FILL
XFILL_15_DFFSR_88 gnd vdd FILL
XFILL_15_DFFSR_99 gnd vdd FILL
XFILL_55_DFFSR_10 gnd vdd FILL
XFILL_55_DFFSR_21 gnd vdd FILL
XFILL_55_DFFSR_32 gnd vdd FILL
XFILL_55_DFFSR_43 gnd vdd FILL
XFILL_26_NOR3X1_7 gnd vdd FILL
XFILL_9_NOR2X1_18 gnd vdd FILL
XFILL_55_DFFSR_54 gnd vdd FILL
XFILL_9_NOR2X1_29 gnd vdd FILL
XFILL_55_DFFSR_65 gnd vdd FILL
XFILL_55_DFFSR_76 gnd vdd FILL
XFILL_55_DFFSR_87 gnd vdd FILL
XFILL_55_DFFSR_98 gnd vdd FILL
XFILL_2_MUX2X1_104 gnd vdd FILL
XFILL_2_MUX2X1_115 gnd vdd FILL
XFILL_44_DFFSR_3 gnd vdd FILL
XFILL_0_NOR2X1_8 gnd vdd FILL
XFILL_2_MUX2X1_126 gnd vdd FILL
XFILL_24_DFFSR_20 gnd vdd FILL
XFILL_2_MUX2X1_137 gnd vdd FILL
XFILL_2_MUX2X1_148 gnd vdd FILL
XFILL_24_DFFSR_31 gnd vdd FILL
XFILL_2_MUX2X1_159 gnd vdd FILL
XFILL_24_DFFSR_42 gnd vdd FILL
XFILL_24_DFFSR_53 gnd vdd FILL
XFILL_24_DFFSR_64 gnd vdd FILL
XFILL_24_DFFSR_75 gnd vdd FILL
XFILL_80_DFFSR_180 gnd vdd FILL
XFILL_24_DFFSR_86 gnd vdd FILL
XFILL_3_OAI21X1_20 gnd vdd FILL
XFILL_80_DFFSR_191 gnd vdd FILL
XFILL_3_OAI21X1_31 gnd vdd FILL
XFILL_31_DFFSR_204 gnd vdd FILL
XFILL_24_DFFSR_97 gnd vdd FILL
XFILL_9_NOR3X1_8 gnd vdd FILL
XFILL_56_3_2 gnd vdd FILL
XFILL_3_OAI21X1_42 gnd vdd FILL
XFILL_31_DFFSR_215 gnd vdd FILL
XFILL_64_DFFSR_30 gnd vdd FILL
XFILL_7_BUFX2_8 gnd vdd FILL
XFILL_31_DFFSR_226 gnd vdd FILL
XFILL_64_DFFSR_41 gnd vdd FILL
XFILL_31_DFFSR_237 gnd vdd FILL
XFILL_0_DFFSR_250 gnd vdd FILL
XFILL_31_DFFSR_248 gnd vdd FILL
XFILL_64_DFFSR_52 gnd vdd FILL
XFILL_0_DFFSR_261 gnd vdd FILL
XFILL_64_DFFSR_63 gnd vdd FILL
XFILL_31_DFFSR_259 gnd vdd FILL
XFILL_0_DFFSR_272 gnd vdd FILL
XFILL_64_DFFSR_74 gnd vdd FILL
XFILL_64_DFFSR_85 gnd vdd FILL
XFILL_84_DFFSR_190 gnd vdd FILL
XFILL_64_DFFSR_96 gnd vdd FILL
XFILL_0_7_0 gnd vdd FILL
XFILL_35_DFFSR_203 gnd vdd FILL
XFILL_25_7_0 gnd vdd FILL
XFILL_35_DFFSR_214 gnd vdd FILL
XFILL_7_DFFSR_10 gnd vdd FILL
XFILL_7_DFFSR_21 gnd vdd FILL
XFILL_35_DFFSR_225 gnd vdd FILL
XFILL_35_DFFSR_236 gnd vdd FILL
XFILL_7_DFFSR_32 gnd vdd FILL
XFILL_35_DFFSR_247 gnd vdd FILL
XFILL_4_DFFSR_260 gnd vdd FILL
XFILL_4_DFFSR_271 gnd vdd FILL
XFILL_7_DFFSR_43 gnd vdd FILL
XFILL_35_DFFSR_258 gnd vdd FILL
XFILL_66_DFFSR_7 gnd vdd FILL
XFILL_35_DFFSR_269 gnd vdd FILL
XFILL_7_DFFSR_54 gnd vdd FILL
XFILL_33_DFFSR_40 gnd vdd FILL
XFILL_7_DFFSR_65 gnd vdd FILL
XFILL_1_MUX2X1_16 gnd vdd FILL
XFILL_7_DFFSR_76 gnd vdd FILL
XFILL_33_DFFSR_51 gnd vdd FILL
XFILL_1_MUX2X1_27 gnd vdd FILL
XFILL_39_DFFSR_202 gnd vdd FILL
XFILL_62_DFFSR_103 gnd vdd FILL
XFILL_7_DFFSR_87 gnd vdd FILL
XFILL_1_MUX2X1_38 gnd vdd FILL
XFILL_39_DFFSR_213 gnd vdd FILL
XFILL_62_DFFSR_114 gnd vdd FILL
XFILL_33_DFFSR_62 gnd vdd FILL
XFILL_7_DFFSR_98 gnd vdd FILL
XFILL_33_DFFSR_73 gnd vdd FILL
XFILL_1_MUX2X1_49 gnd vdd FILL
XFILL_39_DFFSR_224 gnd vdd FILL
XFILL_62_DFFSR_125 gnd vdd FILL
XFILL_62_DFFSR_136 gnd vdd FILL
XFILL_33_DFFSR_84 gnd vdd FILL
XFILL_33_DFFSR_95 gnd vdd FILL
XFILL_39_DFFSR_235 gnd vdd FILL
XFILL_62_DFFSR_147 gnd vdd FILL
XFILL_39_DFFSR_246 gnd vdd FILL
XFILL_62_DFFSR_158 gnd vdd FILL
XFILL_8_DFFSR_270 gnd vdd FILL
XFILL_39_DFFSR_257 gnd vdd FILL
XFILL_39_DFFSR_268 gnd vdd FILL
XFILL_62_DFFSR_169 gnd vdd FILL
XFILL_5_MUX2X1_15 gnd vdd FILL
XFILL_66_DFFSR_102 gnd vdd FILL
XFILL_5_MUX2X1_26 gnd vdd FILL
XFILL_73_DFFSR_50 gnd vdd FILL
XFILL_5_MUX2X1_37 gnd vdd FILL
XFILL_73_DFFSR_61 gnd vdd FILL
XFILL_5_MUX2X1_48 gnd vdd FILL
XFILL_66_DFFSR_113 gnd vdd FILL
XFILL_66_DFFSR_124 gnd vdd FILL
XFILL_5_NAND3X1_18 gnd vdd FILL
XFILL_73_DFFSR_72 gnd vdd FILL
XFILL_73_DFFSR_83 gnd vdd FILL
XFILL_66_DFFSR_135 gnd vdd FILL
XFILL_5_MUX2X1_59 gnd vdd FILL
XFILL_5_NAND3X1_29 gnd vdd FILL
XFILL_66_DFFSR_146 gnd vdd FILL
XFILL_73_DFFSR_94 gnd vdd FILL
XFILL_66_DFFSR_157 gnd vdd FILL
XFILL_66_DFFSR_168 gnd vdd FILL
XFILL_66_DFFSR_179 gnd vdd FILL
XFILL_9_MUX2X1_14 gnd vdd FILL
XFILL_9_MUX2X1_25 gnd vdd FILL
XFILL_6_BUFX4_2 gnd vdd FILL
XFILL_9_MUX2X1_36 gnd vdd FILL
XFILL_9_MUX2X1_47 gnd vdd FILL
XFILL_13_NOR3X1_2 gnd vdd FILL
XFILL_9_MUX2X1_58 gnd vdd FILL
XFILL_13_OAI21X1_2 gnd vdd FILL
XFILL_9_MUX2X1_69 gnd vdd FILL
XFILL_42_DFFSR_60 gnd vdd FILL
XFILL_19_MUX2X1_140 gnd vdd FILL
XFILL_42_DFFSR_71 gnd vdd FILL
XFILL_19_MUX2X1_151 gnd vdd FILL
XFILL_42_DFFSR_82 gnd vdd FILL
XFILL_10_NOR2X1_60 gnd vdd FILL
XFILL_19_MUX2X1_162 gnd vdd FILL
XFILL_42_DFFSR_93 gnd vdd FILL
XFILL_10_NOR2X1_71 gnd vdd FILL
XFILL_19_MUX2X1_173 gnd vdd FILL
XBUFX4_15 BUFX4_54/A gnd DFFSR_26/R vdd BUFX4
XFILL_10_NOR2X1_82 gnd vdd FILL
XFILL_10_NOR2X1_93 gnd vdd FILL
XBUFX4_26 BUFX4_47/A gnd DFFSR_87/R vdd BUFX4
XFILL_19_MUX2X1_184 gnd vdd FILL
XFILL_1_INVX1_220 gnd vdd FILL
XBUFX4_37 BUFX4_44/A gnd DFFSR_1/R vdd BUFX4
XBUFX4_48 BUFX4_54/A gnd DFFSR_25/R vdd BUFX4
XBUFX4_59 BUFX4_60/A gnd INVX2_2/A vdd BUFX4
XFILL_82_DFFSR_70 gnd vdd FILL
XFILL_47_3_2 gnd vdd FILL
XFILL_82_DFFSR_81 gnd vdd FILL
XFILL_82_DFFSR_92 gnd vdd FILL
XFILL_21_MUX2X1_13 gnd vdd FILL
XFILL_5_INVX1_6 gnd vdd FILL
XFILL_11_DFFSR_70 gnd vdd FILL
XFILL_21_MUX2X1_24 gnd vdd FILL
XFILL_21_MUX2X1_35 gnd vdd FILL
XFILL_11_DFFSR_81 gnd vdd FILL
XFILL_21_MUX2X1_46 gnd vdd FILL
XFILL_11_DFFSR_92 gnd vdd FILL
XFILL_21_MUX2X1_57 gnd vdd FILL
XFILL_21_MUX2X1_68 gnd vdd FILL
XFILL_16_7_0 gnd vdd FILL
XFILL_21_MUX2X1_79 gnd vdd FILL
XFILL_51_DFFSR_190 gnd vdd FILL
XFILL_51_DFFSR_80 gnd vdd FILL
XFILL_51_DFFSR_91 gnd vdd FILL
XFILL_30_2_2 gnd vdd FILL
XFILL_24_CLKBUF1_19 gnd vdd FILL
XFILL_20_DFFSR_90 gnd vdd FILL
XFILL_5_NOR3X1_1 gnd vdd FILL
XFILL_9_MUX2X1_190 gnd vdd FILL
XFILL_33_DFFSR_102 gnd vdd FILL
XFILL_10_NAND2X1_4 gnd vdd FILL
XFILL_33_DFFSR_113 gnd vdd FILL
XFILL_33_DFFSR_124 gnd vdd FILL
XFILL_33_DFFSR_135 gnd vdd FILL
XFILL_33_DFFSR_146 gnd vdd FILL
XFILL_33_DFFSR_157 gnd vdd FILL
XFILL_2_DFFSR_170 gnd vdd FILL
XFILL_33_DFFSR_168 gnd vdd FILL
XFILL_2_DFFSR_181 gnd vdd FILL
XFILL_33_DFFSR_179 gnd vdd FILL
XFILL_2_DFFSR_192 gnd vdd FILL
XFILL_37_DFFSR_101 gnd vdd FILL
XFILL_37_DFFSR_112 gnd vdd FILL
XFILL_5_NOR2X1_108 gnd vdd FILL
XFILL_37_DFFSR_123 gnd vdd FILL
XFILL_37_DFFSR_134 gnd vdd FILL
XFILL_5_NOR2X1_119 gnd vdd FILL
XFILL_37_DFFSR_145 gnd vdd FILL
XFILL_11_NAND3X1_10 gnd vdd FILL
XFILL_37_DFFSR_156 gnd vdd FILL
XFILL_11_NAND3X1_21 gnd vdd FILL
XFILL_83_DFFSR_1 gnd vdd FILL
XFILL_6_DFFSR_180 gnd vdd FILL
XFILL_37_DFFSR_167 gnd vdd FILL
XFILL_11_NAND3X1_32 gnd vdd FILL
XFILL_3_DFFSR_80 gnd vdd FILL
XFILL_37_DFFSR_178 gnd vdd FILL
XFILL_6_DFFSR_191 gnd vdd FILL
XFILL_11_NAND3X1_43 gnd vdd FILL
XFILL_3_DFFSR_91 gnd vdd FILL
XFILL_37_DFFSR_189 gnd vdd FILL
XFILL_11_NAND3X1_54 gnd vdd FILL
XFILL_11_NAND3X1_65 gnd vdd FILL
XFILL_31_CLKBUF1_10 gnd vdd FILL
XFILL_66_6_0 gnd vdd FILL
XFILL_11_NAND3X1_76 gnd vdd FILL
XFILL_31_CLKBUF1_21 gnd vdd FILL
XFILL_38_3_2 gnd vdd FILL
XFILL_31_CLKBUF1_32 gnd vdd FILL
XFILL_11_NAND3X1_87 gnd vdd FILL
XFILL_11_NAND3X1_98 gnd vdd FILL
XFILL_83_DFFSR_202 gnd vdd FILL
XFILL_83_DFFSR_213 gnd vdd FILL
XFILL_10_DFFSR_6 gnd vdd FILL
XFILL_83_DFFSR_224 gnd vdd FILL
XFILL_83_DFFSR_235 gnd vdd FILL
XFILL_10_AOI21X1_9 gnd vdd FILL
XFILL_83_DFFSR_246 gnd vdd FILL
XFILL_83_DFFSR_257 gnd vdd FILL
XFILL_83_DFFSR_268 gnd vdd FILL
XFILL_48_DFFSR_4 gnd vdd FILL
XFILL_87_DFFSR_201 gnd vdd FILL
XFILL_87_DFFSR_212 gnd vdd FILL
XFILL_21_2_2 gnd vdd FILL
XFILL_87_DFFSR_223 gnd vdd FILL
XFILL_2_OAI22X1_17 gnd vdd FILL
XFILL_14_AOI21X1_8 gnd vdd FILL
XFILL_87_DFFSR_234 gnd vdd FILL
XFILL_87_DFFSR_245 gnd vdd FILL
XFILL_2_OAI22X1_28 gnd vdd FILL
XFILL_87_DFFSR_256 gnd vdd FILL
XFILL_2_OAI22X1_39 gnd vdd FILL
XFILL_87_DFFSR_267 gnd vdd FILL
XFILL_15_AOI22X1_10 gnd vdd FILL
XFILL_6_OAI21X1_19 gnd vdd FILL
XFILL_3_INVX1_140 gnd vdd FILL
XFILL_3_INVX1_151 gnd vdd FILL
XFILL_3_INVX1_162 gnd vdd FILL
XFILL_3_INVX1_173 gnd vdd FILL
XFILL_1_NAND3X1_60 gnd vdd FILL
XFILL_3_INVX1_184 gnd vdd FILL
XFILL_1_NAND3X1_71 gnd vdd FILL
XFILL_3_INVX1_195 gnd vdd FILL
XFILL_1_NAND3X1_82 gnd vdd FILL
XFILL_1_NAND3X1_93 gnd vdd FILL
XFILL_5_NAND2X1_40 gnd vdd FILL
XFILL_5_NAND2X1_51 gnd vdd FILL
XFILL_5_NAND2X1_62 gnd vdd FILL
XFILL_7_INVX1_150 gnd vdd FILL
XFILL_5_NAND2X1_73 gnd vdd FILL
XFILL_7_INVX1_161 gnd vdd FILL
XFILL_5_NAND2X1_84 gnd vdd FILL
XFILL_5_NAND2X1_95 gnd vdd FILL
XFILL_7_INVX1_172 gnd vdd FILL
XFILL_7_INVX1_183 gnd vdd FILL
XFILL_7_INVX1_194 gnd vdd FILL
XFILL_13_CLKBUF1_15 gnd vdd FILL
XFILL_13_CLKBUF1_26 gnd vdd FILL
XFILL_13_CLKBUF1_37 gnd vdd FILL
XFILL_1_OAI22X1_2 gnd vdd FILL
XFILL_57_6_0 gnd vdd FILL
XFILL_4_3_2 gnd vdd FILL
XFILL_29_3_2 gnd vdd FILL
XFILL_5_OAI22X1_1 gnd vdd FILL
XFILL_11_NOR2X1_100 gnd vdd FILL
XFILL_11_NOR2X1_111 gnd vdd FILL
XFILL_11_NOR2X1_122 gnd vdd FILL
XFILL_11_NOR2X1_133 gnd vdd FILL
XFILL_11_NOR2X1_144 gnd vdd FILL
XFILL_11_NOR2X1_155 gnd vdd FILL
XFILL_11_NOR2X1_166 gnd vdd FILL
XFILL_50_DFFSR_202 gnd vdd FILL
XFILL_11_NOR2X1_177 gnd vdd FILL
XFILL_50_DFFSR_213 gnd vdd FILL
XFILL_11_NOR2X1_188 gnd vdd FILL
XFILL_11_NOR2X1_199 gnd vdd FILL
XFILL_50_DFFSR_224 gnd vdd FILL
XFILL_50_DFFSR_235 gnd vdd FILL
XFILL_40_5_0 gnd vdd FILL
XFILL_9_AOI21X1_40 gnd vdd FILL
XFILL_50_DFFSR_246 gnd vdd FILL
XFILL_65_DFFSR_19 gnd vdd FILL
XFILL_9_AOI21X1_51 gnd vdd FILL
XFILL_12_2_2 gnd vdd FILL
XFILL_50_DFFSR_257 gnd vdd FILL
XFILL_9_AOI21X1_62 gnd vdd FILL
XFILL_50_DFFSR_268 gnd vdd FILL
XFILL_9_AOI21X1_73 gnd vdd FILL
XFILL_19_OAI22X1_20 gnd vdd FILL
XFILL_19_OAI22X1_31 gnd vdd FILL
XFILL_54_DFFSR_201 gnd vdd FILL
XFILL_19_OAI22X1_42 gnd vdd FILL
XFILL_54_DFFSR_212 gnd vdd FILL
XFILL_54_DFFSR_223 gnd vdd FILL
XFILL_54_DFFSR_234 gnd vdd FILL
XFILL_54_DFFSR_245 gnd vdd FILL
XFILL_3_CLKBUF1_10 gnd vdd FILL
XFILL_54_DFFSR_256 gnd vdd FILL
XFILL_3_CLKBUF1_21 gnd vdd FILL
XFILL_54_DFFSR_267 gnd vdd FILL
XFILL_3_CLKBUF1_32 gnd vdd FILL
XFILL_81_DFFSR_101 gnd vdd FILL
XFILL_58_DFFSR_200 gnd vdd FILL
XFILL_58_DFFSR_211 gnd vdd FILL
XFILL_11_MUX2X1_106 gnd vdd FILL
XFILL_34_DFFSR_18 gnd vdd FILL
XFILL_81_DFFSR_112 gnd vdd FILL
XFILL_11_MUX2X1_117 gnd vdd FILL
XFILL_58_DFFSR_222 gnd vdd FILL
XFILL_34_DFFSR_29 gnd vdd FILL
XFILL_81_DFFSR_123 gnd vdd FILL
XFILL_81_DFFSR_134 gnd vdd FILL
XFILL_11_MUX2X1_128 gnd vdd FILL
XFILL_58_DFFSR_233 gnd vdd FILL
XFILL_81_DFFSR_145 gnd vdd FILL
XFILL_11_MUX2X1_139 gnd vdd FILL
XFILL_58_DFFSR_244 gnd vdd FILL
XFILL_81_DFFSR_156 gnd vdd FILL
XFILL_58_DFFSR_255 gnd vdd FILL
XFILL_81_DFFSR_167 gnd vdd FILL
XFILL_58_DFFSR_266 gnd vdd FILL
XFILL_13_CLKBUF1_7 gnd vdd FILL
XFILL_81_DFFSR_178 gnd vdd FILL
XFILL_85_DFFSR_100 gnd vdd FILL
XFILL_81_DFFSR_189 gnd vdd FILL
XFILL_1_DFFSR_204 gnd vdd FILL
XFILL_1_DFFSR_215 gnd vdd FILL
XFILL_12_OAI21X1_11 gnd vdd FILL
XFILL_74_DFFSR_17 gnd vdd FILL
XFILL_85_DFFSR_111 gnd vdd FILL
XFILL_74_DFFSR_28 gnd vdd FILL
XFILL_1_DFFSR_226 gnd vdd FILL
XFILL_85_DFFSR_122 gnd vdd FILL
XFILL_12_OAI21X1_22 gnd vdd FILL
XFILL_85_DFFSR_133 gnd vdd FILL
XFILL_1_DFFSR_237 gnd vdd FILL
XFILL_74_DFFSR_39 gnd vdd FILL
XFILL_12_OAI21X1_33 gnd vdd FILL
XFILL_85_DFFSR_144 gnd vdd FILL
XFILL_1_DFFSR_248 gnd vdd FILL
XFILL_85_DFFSR_155 gnd vdd FILL
XFILL_1_NOR2X1_150 gnd vdd FILL
XFILL_12_OAI21X1_44 gnd vdd FILL
XFILL_1_DFFSR_259 gnd vdd FILL
XFILL_17_MUX2X1_7 gnd vdd FILL
XFILL_1_NOR2X1_161 gnd vdd FILL
XFILL_85_DFFSR_166 gnd vdd FILL
XFILL_85_DFFSR_177 gnd vdd FILL
XFILL_1_NOR2X1_172 gnd vdd FILL
XFILL_17_CLKBUF1_6 gnd vdd FILL
XFILL_1_NOR2X1_183 gnd vdd FILL
XFILL_85_DFFSR_188 gnd vdd FILL
XFILL_5_DFFSR_203 gnd vdd FILL
XFILL_2_NAND3X1_3 gnd vdd FILL
XFILL_1_NOR2X1_194 gnd vdd FILL
XFILL_85_DFFSR_199 gnd vdd FILL
XFILL_5_DFFSR_214 gnd vdd FILL
XFILL_48_6_0 gnd vdd FILL
XFILL_5_DFFSR_225 gnd vdd FILL
XFILL_8_BUFX4_40 gnd vdd FILL
XFILL_5_DFFSR_236 gnd vdd FILL
XFILL_8_BUFX4_51 gnd vdd FILL
XFILL_5_DFFSR_247 gnd vdd FILL
XFILL_13_BUFX4_101 gnd vdd FILL
XFILL_5_DFFSR_258 gnd vdd FILL
XFILL_8_BUFX4_62 gnd vdd FILL
XFILL_5_DFFSR_269 gnd vdd FILL
XFILL_8_BUFX4_73 gnd vdd FILL
XFILL_43_DFFSR_16 gnd vdd FILL
XFILL_43_DFFSR_27 gnd vdd FILL
XFILL_8_BUFX4_84 gnd vdd FILL
XFILL_43_DFFSR_38 gnd vdd FILL
XFILL_9_DFFSR_202 gnd vdd FILL
XFILL_8_BUFX4_95 gnd vdd FILL
XFILL_43_DFFSR_49 gnd vdd FILL
XFILL_9_DFFSR_213 gnd vdd FILL
XFILL_6_NAND3X1_2 gnd vdd FILL
XFILL_9_DFFSR_224 gnd vdd FILL
XFILL_62_1_2 gnd vdd FILL
XFILL_9_DFFSR_235 gnd vdd FILL
XFILL_9_DFFSR_246 gnd vdd FILL
XFILL_83_DFFSR_15 gnd vdd FILL
XFILL_9_DFFSR_257 gnd vdd FILL
XFILL_9_DFFSR_268 gnd vdd FILL
XFILL_83_DFFSR_26 gnd vdd FILL
XFILL_83_DFFSR_37 gnd vdd FILL
XFILL_1_MUX2X1_101 gnd vdd FILL
XFILL_1_MUX2X1_112 gnd vdd FILL
XFILL_83_DFFSR_48 gnd vdd FILL
XFILL_1_MUX2X1_123 gnd vdd FILL
XFILL_12_DFFSR_15 gnd vdd FILL
XFILL_83_DFFSR_59 gnd vdd FILL
XFILL_31_5_0 gnd vdd FILL
XFILL_12_DFFSR_26 gnd vdd FILL
XFILL_1_MUX2X1_134 gnd vdd FILL
XFILL_1_MUX2X1_145 gnd vdd FILL
XFILL_12_DFFSR_37 gnd vdd FILL
XFILL_1_MUX2X1_156 gnd vdd FILL
XFILL_12_DFFSR_48 gnd vdd FILL
XFILL_1_MUX2X1_167 gnd vdd FILL
XFILL_87_DFFSR_2 gnd vdd FILL
XFILL_12_DFFSR_59 gnd vdd FILL
XFILL_1_MUX2X1_178 gnd vdd FILL
XFILL_1_MUX2X1_189 gnd vdd FILL
XFILL_52_DFFSR_14 gnd vdd FILL
XFILL_21_DFFSR_201 gnd vdd FILL
XFILL_52_DFFSR_25 gnd vdd FILL
XFILL_21_DFFSR_212 gnd vdd FILL
XFILL_2_OAI21X1_50 gnd vdd FILL
XFILL_52_DFFSR_36 gnd vdd FILL
XFILL_11_NOR2X1_14 gnd vdd FILL
XFILL_11_NOR2X1_25 gnd vdd FILL
XFILL_21_DFFSR_223 gnd vdd FILL
XFILL_2_AOI22X1_8 gnd vdd FILL
XFILL_52_DFFSR_47 gnd vdd FILL
XFILL_21_DFFSR_234 gnd vdd FILL
XFILL_52_DFFSR_58 gnd vdd FILL
XFILL_11_NOR2X1_36 gnd vdd FILL
XFILL_11_NOR2X1_47 gnd vdd FILL
XFILL_52_DFFSR_69 gnd vdd FILL
XFILL_21_DFFSR_245 gnd vdd FILL
XFILL_21_DFFSR_256 gnd vdd FILL
XFILL_11_NOR2X1_58 gnd vdd FILL
XFILL_21_DFFSR_267 gnd vdd FILL
XFILL_11_NOR2X1_69 gnd vdd FILL
XFILL_2_INVX1_207 gnd vdd FILL
XFILL_25_DFFSR_200 gnd vdd FILL
XFILL_25_DFFSR_211 gnd vdd FILL
XFILL_1_DFFSR_9 gnd vdd FILL
XFILL_9_MUX2X1_6 gnd vdd FILL
XFILL_2_INVX1_218 gnd vdd FILL
XFILL_25_DFFSR_222 gnd vdd FILL
XFILL_14_DFFSR_7 gnd vdd FILL
XFILL_6_AOI22X1_7 gnd vdd FILL
XFILL_21_DFFSR_13 gnd vdd FILL
XFILL_25_DFFSR_233 gnd vdd FILL
XFILL_21_DFFSR_24 gnd vdd FILL
XFILL_71_DFFSR_8 gnd vdd FILL
XFILL_25_DFFSR_244 gnd vdd FILL
XFILL_21_DFFSR_35 gnd vdd FILL
XFILL_25_DFFSR_255 gnd vdd FILL
XFILL_25_DFFSR_266 gnd vdd FILL
XFILL_21_DFFSR_46 gnd vdd FILL
XFILL_6_INVX1_206 gnd vdd FILL
XFILL_21_DFFSR_57 gnd vdd FILL
XFILL_52_DFFSR_100 gnd vdd FILL
XFILL_21_DFFSR_68 gnd vdd FILL
XFILL_6_INVX1_217 gnd vdd FILL
XFILL_29_DFFSR_210 gnd vdd FILL
XFILL_52_DFFSR_111 gnd vdd FILL
XFILL_21_DFFSR_79 gnd vdd FILL
XFILL_29_DFFSR_221 gnd vdd FILL
XFILL_6_INVX1_228 gnd vdd FILL
XFILL_52_DFFSR_122 gnd vdd FILL
XFILL_52_DFFSR_133 gnd vdd FILL
XFILL_29_DFFSR_232 gnd vdd FILL
XFILL_52_DFFSR_144 gnd vdd FILL
XFILL_61_DFFSR_12 gnd vdd FILL
XFILL_29_DFFSR_243 gnd vdd FILL
XFILL_61_DFFSR_23 gnd vdd FILL
XFILL_52_DFFSR_155 gnd vdd FILL
XFILL_29_DFFSR_254 gnd vdd FILL
XFILL_39_6_0 gnd vdd FILL
XFILL_61_DFFSR_34 gnd vdd FILL
XFILL_61_DFFSR_45 gnd vdd FILL
XFILL_52_DFFSR_166 gnd vdd FILL
XFILL_29_DFFSR_265 gnd vdd FILL
XFILL_52_DFFSR_177 gnd vdd FILL
XFILL_61_DFFSR_56 gnd vdd FILL
XFILL_52_DFFSR_188 gnd vdd FILL
XFILL_61_DFFSR_67 gnd vdd FILL
XFILL_56_DFFSR_110 gnd vdd FILL
XFILL_52_DFFSR_199 gnd vdd FILL
XFILL_61_DFFSR_78 gnd vdd FILL
XFILL_61_DFFSR_89 gnd vdd FILL
XFILL_4_NAND3X1_15 gnd vdd FILL
XFILL_56_DFFSR_121 gnd vdd FILL
XFILL_56_DFFSR_132 gnd vdd FILL
XFILL_4_NAND3X1_26 gnd vdd FILL
XFILL_56_DFFSR_143 gnd vdd FILL
XFILL_4_NAND3X1_37 gnd vdd FILL
XFILL_56_DFFSR_154 gnd vdd FILL
XFILL_4_DFFSR_14 gnd vdd FILL
XFILL_4_NAND3X1_48 gnd vdd FILL
XFILL_53_1_2 gnd vdd FILL
XFILL_4_NAND3X1_59 gnd vdd FILL
XFILL_56_DFFSR_165 gnd vdd FILL
XFILL_4_DFFSR_25 gnd vdd FILL
XFILL_8_NAND2X1_17 gnd vdd FILL
XFILL_4_DFFSR_36 gnd vdd FILL
XFILL_56_DFFSR_176 gnd vdd FILL
XFILL_8_NAND2X1_28 gnd vdd FILL
XFILL_30_DFFSR_11 gnd vdd FILL
XFILL_56_DFFSR_187 gnd vdd FILL
XFILL_56_DFFSR_198 gnd vdd FILL
XFILL_30_DFFSR_22 gnd vdd FILL
XFILL_8_NAND2X1_39 gnd vdd FILL
XFILL_4_DFFSR_47 gnd vdd FILL
XFILL_4_DFFSR_58 gnd vdd FILL
XFILL_30_DFFSR_33 gnd vdd FILL
XFILL_4_DFFSR_69 gnd vdd FILL
XFILL_30_DFFSR_44 gnd vdd FILL
XFILL_30_DFFSR_55 gnd vdd FILL
XFILL_30_DFFSR_66 gnd vdd FILL
XFILL_30_DFFSR_77 gnd vdd FILL
XFILL_22_5_0 gnd vdd FILL
XFILL_30_DFFSR_88 gnd vdd FILL
XFILL_3_DFFSR_102 gnd vdd FILL
XFILL_30_DFFSR_99 gnd vdd FILL
XFILL_6_INVX1_90 gnd vdd FILL
XFILL_70_DFFSR_10 gnd vdd FILL
XFILL_6_BUFX2_10 gnd vdd FILL
XFILL_70_DFFSR_21 gnd vdd FILL
XFILL_18_MUX2X1_170 gnd vdd FILL
XFILL_3_DFFSR_113 gnd vdd FILL
XFILL_3_DFFSR_124 gnd vdd FILL
XFILL_70_DFFSR_32 gnd vdd FILL
XFILL_18_MUX2X1_181 gnd vdd FILL
XFILL_70_DFFSR_43 gnd vdd FILL
XFILL_3_DFFSR_135 gnd vdd FILL
XFILL_18_MUX2X1_192 gnd vdd FILL
XFILL_3_DFFSR_146 gnd vdd FILL
XFILL_70_DFFSR_54 gnd vdd FILL
XFILL_70_DFFSR_65 gnd vdd FILL
XFILL_3_DFFSR_157 gnd vdd FILL
XFILL_70_DFFSR_76 gnd vdd FILL
XFILL_3_DFFSR_168 gnd vdd FILL
XFILL_3_DFFSR_179 gnd vdd FILL
XFILL_70_DFFSR_87 gnd vdd FILL
XFILL_70_DFFSR_98 gnd vdd FILL
XFILL_7_DFFSR_101 gnd vdd FILL
XFILL_11_MUX2X1_10 gnd vdd FILL
XFILL_7_DFFSR_112 gnd vdd FILL
XFILL_11_MUX2X1_21 gnd vdd FILL
XFILL_7_DFFSR_123 gnd vdd FILL
XFILL_7_DFFSR_134 gnd vdd FILL
XFILL_11_MUX2X1_32 gnd vdd FILL
XFILL_7_DFFSR_145 gnd vdd FILL
XFILL_11_MUX2X1_43 gnd vdd FILL
XFILL_7_DFFSR_156 gnd vdd FILL
XDFFSR_170 INVX1_46/A DFFSR_56/CLK DFFSR_56/R vdd MUX2X1_13/Y gnd vdd DFFSR
XFILL_11_MUX2X1_54 gnd vdd FILL
XFILL_7_DFFSR_167 gnd vdd FILL
XFILL_11_MUX2X1_65 gnd vdd FILL
XDFFSR_181 DFFSR_181/Q DFFSR_58/CLK DFFSR_55/R vdd DFFSR_181/D gnd vdd DFFSR
XFILL_7_DFFSR_178 gnd vdd FILL
XFILL_11_MUX2X1_76 gnd vdd FILL
XFILL_10_NOR3X1_6 gnd vdd FILL
XDFFSR_192 INVX1_131/A DFFSR_90/CLK BUFX4_32/Y vdd DFFSR_192/D gnd vdd DFFSR
XFILL_11_MUX2X1_87 gnd vdd FILL
XFILL_7_DFFSR_189 gnd vdd FILL
XFILL_11_MUX2X1_98 gnd vdd FILL
XFILL_15_MUX2X1_20 gnd vdd FILL
XFILL_15_MUX2X1_31 gnd vdd FILL
XFILL_15_MUX2X1_42 gnd vdd FILL
XFILL_15_MUX2X1_53 gnd vdd FILL
XFILL_15_MUX2X1_64 gnd vdd FILL
XFILL_3_NOR3X1_13 gnd vdd FILL
XFILL_15_MUX2X1_75 gnd vdd FILL
XFILL_15_MUX2X1_86 gnd vdd FILL
XFILL_3_NOR3X1_24 gnd vdd FILL
XFILL_15_MUX2X1_97 gnd vdd FILL
XFILL_3_NOR3X1_35 gnd vdd FILL
XFILL_3_NOR3X1_46 gnd vdd FILL
XFILL_23_CLKBUF1_16 gnd vdd FILL
XFILL_19_MUX2X1_30 gnd vdd FILL
XFILL_5_6_0 gnd vdd FILL
XFILL_19_MUX2X1_41 gnd vdd FILL
XFILL_23_CLKBUF1_27 gnd vdd FILL
XFILL_23_CLKBUF1_38 gnd vdd FILL
XFILL_19_MUX2X1_52 gnd vdd FILL
XFILL_6_NOR2X1_1 gnd vdd FILL
XFILL_19_MUX2X1_63 gnd vdd FILL
XFILL_7_NOR3X1_12 gnd vdd FILL
XFILL_19_MUX2X1_74 gnd vdd FILL
XFILL_19_MUX2X1_85 gnd vdd FILL
XFILL_7_NOR3X1_23 gnd vdd FILL
XFILL_7_NOR3X1_34 gnd vdd FILL
XFILL_19_MUX2X1_96 gnd vdd FILL
XFILL_0_INVX1_106 gnd vdd FILL
XFILL_0_INVX1_117 gnd vdd FILL
XFILL_7_NOR3X1_45 gnd vdd FILL
XFILL_0_INVX1_128 gnd vdd FILL
XFILL_23_DFFSR_110 gnd vdd FILL
XFILL_1_AOI21X1_17 gnd vdd FILL
XFILL_0_INVX1_139 gnd vdd FILL
XFILL_23_DFFSR_121 gnd vdd FILL
XFILL_44_1_2 gnd vdd FILL
XFILL_23_DFFSR_132 gnd vdd FILL
XFILL_23_DFFSR_143 gnd vdd FILL
XFILL_1_AOI21X1_28 gnd vdd FILL
XFILL_23_DFFSR_154 gnd vdd FILL
XFILL_1_AOI21X1_39 gnd vdd FILL
XFILL_23_DFFSR_165 gnd vdd FILL
XFILL_4_INVX1_105 gnd vdd FILL
XFILL_11_OAI22X1_19 gnd vdd FILL
XFILL_23_DFFSR_176 gnd vdd FILL
XFILL_23_DFFSR_187 gnd vdd FILL
XFILL_23_DFFSR_198 gnd vdd FILL
XFILL_4_INVX1_116 gnd vdd FILL
XFILL_4_INVX1_127 gnd vdd FILL
XFILL_4_NOR2X1_105 gnd vdd FILL
XFILL_27_DFFSR_120 gnd vdd FILL
XFILL_13_5_0 gnd vdd FILL
XFILL_4_INVX1_138 gnd vdd FILL
XFILL_27_DFFSR_131 gnd vdd FILL
XFILL_4_NOR2X1_116 gnd vdd FILL
XFILL_31_DFFSR_1 gnd vdd FILL
XFILL_4_INVX1_149 gnd vdd FILL
XFILL_27_DFFSR_142 gnd vdd FILL
XFILL_4_NOR2X1_127 gnd vdd FILL
XFILL_27_DFFSR_153 gnd vdd FILL
XFILL_4_NOR2X1_138 gnd vdd FILL
XFILL_4_NOR2X1_149 gnd vdd FILL
XFILL_27_DFFSR_164 gnd vdd FILL
XFILL_27_DFFSR_175 gnd vdd FILL
XFILL_10_NAND3X1_40 gnd vdd FILL
XFILL_27_DFFSR_186 gnd vdd FILL
XFILL_10_NAND3X1_51 gnd vdd FILL
XFILL_10_NAND3X1_62 gnd vdd FILL
XFILL_27_DFFSR_197 gnd vdd FILL
XFILL_10_NAND3X1_73 gnd vdd FILL
XFILL_2_NOR3X1_5 gnd vdd FILL
XFILL_10_NAND3X1_84 gnd vdd FILL
XFILL_10_NAND3X1_95 gnd vdd FILL
XFILL_30_CLKBUF1_40 gnd vdd FILL
XFILL_23_NOR3X1_10 gnd vdd FILL
XFILL_23_NOR3X1_21 gnd vdd FILL
XFILL_23_NOR3X1_32 gnd vdd FILL
XFILL_23_NOR3X1_43 gnd vdd FILL
XFILL_21_MUX2X1_107 gnd vdd FILL
XFILL_73_DFFSR_210 gnd vdd FILL
XFILL_21_MUX2X1_118 gnd vdd FILL
XFILL_73_DFFSR_221 gnd vdd FILL
XFILL_21_MUX2X1_129 gnd vdd FILL
XFILL_73_DFFSR_232 gnd vdd FILL
XFILL_73_DFFSR_243 gnd vdd FILL
XFILL_0_DFFSR_40 gnd vdd FILL
XFILL_0_DFFSR_51 gnd vdd FILL
XFILL_73_DFFSR_254 gnd vdd FILL
XFILL_73_DFFSR_265 gnd vdd FILL
XFILL_27_NOR3X1_20 gnd vdd FILL
XFILL_53_DFFSR_5 gnd vdd FILL
XFILL_27_NOR3X1_31 gnd vdd FILL
XFILL_0_DFFSR_62 gnd vdd FILL
XFILL_0_DFFSR_73 gnd vdd FILL
XFILL_27_NOR3X1_42 gnd vdd FILL
XFILL_0_DFFSR_84 gnd vdd FILL
XFILL_7_3 gnd vdd FILL
XFILL_0_DFFSR_95 gnd vdd FILL
XFILL_9_NOR2X1_205 gnd vdd FILL
XFILL_77_DFFSR_220 gnd vdd FILL
XFILL_1_OAI22X1_14 gnd vdd FILL
XFILL_77_DFFSR_231 gnd vdd FILL
XFILL_1_OAI22X1_25 gnd vdd FILL
XFILL_63_5 gnd vdd FILL
XFILL_77_DFFSR_242 gnd vdd FILL
XFILL_77_DFFSR_253 gnd vdd FILL
XFILL_1_OAI22X1_36 gnd vdd FILL
XFILL_1_OAI22X1_47 gnd vdd FILL
XFILL_77_DFFSR_264 gnd vdd FILL
XFILL_77_DFFSR_275 gnd vdd FILL
XFILL_32_CLKBUF1_5 gnd vdd FILL
XFILL_5_OAI21X1_16 gnd vdd FILL
XFILL_56_4 gnd vdd FILL
XFILL_5_OAI21X1_27 gnd vdd FILL
XFILL_5_OAI21X1_38 gnd vdd FILL
XFILL_5_OAI21X1_49 gnd vdd FILL
XFILL_63_4_0 gnd vdd FILL
XFILL_35_1_2 gnd vdd FILL
XFILL_0_NAND3X1_90 gnd vdd FILL
XFILL_4_NAND2X1_70 gnd vdd FILL
XFILL_4_NAND2X1_81 gnd vdd FILL
XFILL_18_DFFSR_8 gnd vdd FILL
XFILL_75_DFFSR_9 gnd vdd FILL
XFILL_4_NAND2X1_92 gnd vdd FILL
XFILL_9_BUFX4_18 gnd vdd FILL
XFILL_9_BUFX4_29 gnd vdd FILL
XFILL_12_CLKBUF1_12 gnd vdd FILL
XFILL_12_CLKBUF1_23 gnd vdd FILL
XFILL_59_DFFSR_209 gnd vdd FILL
XFILL_12_CLKBUF1_34 gnd vdd FILL
XFILL_86_DFFSR_109 gnd vdd FILL
XFILL_10_NOR2X1_130 gnd vdd FILL
XFILL_10_NOR2X1_141 gnd vdd FILL
XFILL_10_NOR2X1_152 gnd vdd FILL
XFILL_10_NOR2X1_163 gnd vdd FILL
XFILL_10_NOR2X1_174 gnd vdd FILL
XFILL_40_DFFSR_210 gnd vdd FILL
XFILL_10_NOR2X1_185 gnd vdd FILL
XFILL_10_NOR2X1_196 gnd vdd FILL
XFILL_40_DFFSR_221 gnd vdd FILL
XFILL_40_DFFSR_232 gnd vdd FILL
XFILL_40_DFFSR_243 gnd vdd FILL
XFILL_40_DFFSR_254 gnd vdd FILL
XNAND3X1_3 NAND3X1_3/A BUFX4_2/Y NOR2X1_29/Y gnd NAND3X1_3/Y vdd NAND3X1
XFILL_40_DFFSR_265 gnd vdd FILL
XFILL_8_AOI21X1_70 gnd vdd FILL
XFILL_8_AOI21X1_81 gnd vdd FILL
XFILL_18_OAI22X1_50 gnd vdd FILL
XFILL_44_DFFSR_220 gnd vdd FILL
XFILL_44_DFFSR_231 gnd vdd FILL
XFILL_44_DFFSR_242 gnd vdd FILL
XFILL_44_DFFSR_253 gnd vdd FILL
XFILL_13_BUFX4_12 gnd vdd FILL
XFILL_44_DFFSR_264 gnd vdd FILL
XFILL_44_DFFSR_275 gnd vdd FILL
XFILL_13_BUFX4_23 gnd vdd FILL
XFILL_3_NOR2X1_90 gnd vdd FILL
XFILL_13_BUFX4_34 gnd vdd FILL
XFILL_13_BUFX4_45 gnd vdd FILL
XFILL_10_MUX2X1_103 gnd vdd FILL
XFILL_2_CLKBUF1_40 gnd vdd FILL
XFILL_12_BUFX4_8 gnd vdd FILL
XFILL_54_4_0 gnd vdd FILL
XFILL_13_BUFX4_56 gnd vdd FILL
XFILL_10_MUX2X1_114 gnd vdd FILL
XFILL_71_DFFSR_120 gnd vdd FILL
XFILL_26_1_2 gnd vdd FILL
XFILL_71_DFFSR_131 gnd vdd FILL
XFILL_10_MUX2X1_125 gnd vdd FILL
XFILL_1_1_2 gnd vdd FILL
XFILL_48_DFFSR_230 gnd vdd FILL
XFILL_13_BUFX4_67 gnd vdd FILL
XFILL_71_DFFSR_142 gnd vdd FILL
XFILL_13_BUFX4_78 gnd vdd FILL
XFILL_10_MUX2X1_136 gnd vdd FILL
XFILL_71_DFFSR_153 gnd vdd FILL
XFILL_48_DFFSR_241 gnd vdd FILL
XFILL_13_BUFX4_89 gnd vdd FILL
XFILL_10_MUX2X1_147 gnd vdd FILL
XFILL_10_MUX2X1_158 gnd vdd FILL
XFILL_48_DFFSR_252 gnd vdd FILL
XFILL_48_DFFSR_263 gnd vdd FILL
XFILL_71_DFFSR_164 gnd vdd FILL
XFILL_48_DFFSR_274 gnd vdd FILL
XFILL_71_DFFSR_175 gnd vdd FILL
XFILL_10_MUX2X1_169 gnd vdd FILL
XFILL_71_DFFSR_186 gnd vdd FILL
XFILL_71_DFFSR_197 gnd vdd FILL
XFILL_75_DFFSR_130 gnd vdd FILL
XFILL_11_OAI21X1_30 gnd vdd FILL
XFILL_11_OAI21X1_41 gnd vdd FILL
XFILL_75_DFFSR_141 gnd vdd FILL
XFILL_75_DFFSR_152 gnd vdd FILL
XFILL_75_DFFSR_163 gnd vdd FILL
XFILL_75_DFFSR_174 gnd vdd FILL
XFILL_0_NOR2X1_180 gnd vdd FILL
XFILL_75_DFFSR_185 gnd vdd FILL
XFILL_0_NOR2X1_191 gnd vdd FILL
XFILL_75_DFFSR_196 gnd vdd FILL
XFILL_26_DFFSR_209 gnd vdd FILL
XAOI22X1_8 NOR2X1_40/Y INVX1_178/A INVX1_173/A NOR2X1_41/Y gnd AOI22X1_8/Y vdd AOI22X1
XFILL_79_DFFSR_140 gnd vdd FILL
XFILL_7_INVX1_13 gnd vdd FILL
XFILL_79_DFFSR_151 gnd vdd FILL
XFILL_79_DFFSR_162 gnd vdd FILL
XFILL_7_INVX1_24 gnd vdd FILL
XFILL_7_INVX1_35 gnd vdd FILL
XFILL_79_DFFSR_173 gnd vdd FILL
XINVX1_207 INVX1_207/A gnd OAI22X1_4/C vdd INVX1
XFILL_79_DFFSR_184 gnd vdd FILL
XFILL_7_INVX1_46 gnd vdd FILL
XFILL_8_AND2X2_5 gnd vdd FILL
XINVX1_218 INVX1_218/A gnd INVX1_218/Y vdd INVX1
XFILL_79_DFFSR_195 gnd vdd FILL
XFILL_7_INVX1_57 gnd vdd FILL
XFILL_53_DFFSR_109 gnd vdd FILL
XFILL_7_INVX1_68 gnd vdd FILL
XFILL_7_INVX1_79 gnd vdd FILL
XFILL_9_2_2 gnd vdd FILL
XFILL_0_MUX2X1_120 gnd vdd FILL
XFILL_57_DFFSR_108 gnd vdd FILL
XFILL_3_NAND2X1_1 gnd vdd FILL
XFILL_0_MUX2X1_131 gnd vdd FILL
XFILL_57_DFFSR_119 gnd vdd FILL
XFILL_35_DFFSR_2 gnd vdd FILL
XFILL_5_BUFX4_11 gnd vdd FILL
XFILL_0_MUX2X1_142 gnd vdd FILL
XFILL_0_MUX2X1_153 gnd vdd FILL
XFILL_5_BUFX4_22 gnd vdd FILL
XFILL_0_MUX2X1_164 gnd vdd FILL
XFILL_13_NAND3X1_17 gnd vdd FILL
XNAND2X1_18 NAND3X1_78/Y OAI21X1_34/Y gnd NAND3X1_43/A vdd NAND2X1
XFILL_0_MUX2X1_175 gnd vdd FILL
XFILL_5_BUFX4_33 gnd vdd FILL
XFILL_13_NAND3X1_28 gnd vdd FILL
XFILL_5_BUFX4_44 gnd vdd FILL
XNAND2X1_29 BUFX4_103/Y AND2X2_1/Y gnd OAI22X1_9/D vdd NAND2X1
XFILL_0_MUX2X1_186 gnd vdd FILL
XFILL_13_NAND3X1_39 gnd vdd FILL
XFILL_5_BUFX4_55 gnd vdd FILL
XFILL_5_BUFX4_66 gnd vdd FILL
XFILL_5_BUFX4_77 gnd vdd FILL
XFILL_33_CLKBUF1_17 gnd vdd FILL
XFILL_5_BUFX4_88 gnd vdd FILL
XFILL_33_CLKBUF1_28 gnd vdd FILL
XFILL_5_BUFX4_99 gnd vdd FILL
XFILL_11_DFFSR_220 gnd vdd FILL
XFILL_33_CLKBUF1_39 gnd vdd FILL
XFILL_11_DFFSR_231 gnd vdd FILL
XFILL_11_DFFSR_242 gnd vdd FILL
XFILL_11_DFFSR_253 gnd vdd FILL
XFILL_45_4_0 gnd vdd FILL
XFILL_11_DFFSR_264 gnd vdd FILL
XFILL_80_DFFSR_19 gnd vdd FILL
XFILL_17_1_2 gnd vdd FILL
XFILL_11_DFFSR_275 gnd vdd FILL
XFILL_15_DFFSR_230 gnd vdd FILL
XFILL_23_MUX2X1_9 gnd vdd FILL
XFILL_15_DFFSR_241 gnd vdd FILL
XFILL_15_DFFSR_252 gnd vdd FILL
XFILL_28_8 gnd vdd FILL
XFILL_15_DFFSR_263 gnd vdd FILL
XFILL_15_DFFSR_274 gnd vdd FILL
XFILL_57_DFFSR_6 gnd vdd FILL
XFILL_12_MUX2X1_19 gnd vdd FILL
XFILL_42_DFFSR_130 gnd vdd FILL
XFILL_3_AOI21X1_6 gnd vdd FILL
XFILL_42_DFFSR_141 gnd vdd FILL
XFILL_42_DFFSR_152 gnd vdd FILL
XFILL_19_DFFSR_240 gnd vdd FILL
XFILL_19_DFFSR_251 gnd vdd FILL
XFILL_19_DFFSR_262 gnd vdd FILL
XFILL_42_DFFSR_163 gnd vdd FILL
XFILL_42_DFFSR_174 gnd vdd FILL
XFILL_19_DFFSR_273 gnd vdd FILL
XFILL_42_DFFSR_185 gnd vdd FILL
XFILL_16_MUX2X1_18 gnd vdd FILL
XFILL_42_DFFSR_196 gnd vdd FILL
XFILL_16_MUX2X1_29 gnd vdd FILL
XFILL_3_NAND3X1_12 gnd vdd FILL
XFILL_7_AOI21X1_5 gnd vdd FILL
XFILL_3_NAND3X1_23 gnd vdd FILL
XFILL_46_DFFSR_140 gnd vdd FILL
XFILL_3_NAND3X1_34 gnd vdd FILL
XFILL_46_DFFSR_151 gnd vdd FILL
XNOR3X1_6 NOR3X1_6/A NOR3X1_6/B NOR3X1_6/C gnd NOR3X1_7/C vdd NOR3X1
XFILL_3_NAND3X1_45 gnd vdd FILL
XFILL_46_DFFSR_162 gnd vdd FILL
XFILL_7_NAND2X1_14 gnd vdd FILL
XFILL_3_NAND3X1_56 gnd vdd FILL
XFILL_46_DFFSR_173 gnd vdd FILL
XFILL_3_NAND3X1_67 gnd vdd FILL
XFILL_7_NAND2X1_25 gnd vdd FILL
XFILL_46_DFFSR_184 gnd vdd FILL
XFILL_3_NAND3X1_78 gnd vdd FILL
XFILL_3_NAND3X1_89 gnd vdd FILL
XFILL_46_DFFSR_195 gnd vdd FILL
XFILL_7_NAND2X1_36 gnd vdd FILL
XFILL_20_DFFSR_109 gnd vdd FILL
XFILL_7_NAND2X1_47 gnd vdd FILL
XFILL_7_NAND2X1_58 gnd vdd FILL
XFILL_7_NAND2X1_69 gnd vdd FILL
XFILL_12_AOI22X1_2 gnd vdd FILL
XFILL_24_DFFSR_108 gnd vdd FILL
XFILL_24_DFFSR_119 gnd vdd FILL
XFILL_61_2 gnd vdd FILL
XFILL_16_AOI22X1_1 gnd vdd FILL
XFILL_10_AOI21X1_19 gnd vdd FILL
XFILL_54_1 gnd vdd FILL
XFILL_28_DFFSR_107 gnd vdd FILL
XFILL_1_DFFSR_18 gnd vdd FILL
XFILL_1_DFFSR_29 gnd vdd FILL
XFILL_11_NOR2X1_6 gnd vdd FILL
XFILL_28_DFFSR_118 gnd vdd FILL
XFILL_36_4_0 gnd vdd FILL
XFILL_28_DFFSR_129 gnd vdd FILL
XFILL_3_INVX1_50 gnd vdd FILL
XFILL_3_INVX1_61 gnd vdd FILL
XFILL_3_INVX1_72 gnd vdd FILL
XFILL_3_INVX1_83 gnd vdd FILL
XFILL_49_DFFSR_20 gnd vdd FILL
XFILL_3_INVX1_94 gnd vdd FILL
XFILL_49_DFFSR_31 gnd vdd FILL
XFILL_70_DFFSR_209 gnd vdd FILL
XFILL_49_DFFSR_42 gnd vdd FILL
XFILL_49_DFFSR_53 gnd vdd FILL
XFILL_49_DFFSR_64 gnd vdd FILL
XFILL_10_MUX2X1_4 gnd vdd FILL
XFILL_49_DFFSR_75 gnd vdd FILL
XFILL_49_DFFSR_86 gnd vdd FILL
XFILL_24_NOR3X1_19 gnd vdd FILL
XFILL_49_DFFSR_97 gnd vdd FILL
XFILL_22_CLKBUF1_13 gnd vdd FILL
XFILL_74_DFFSR_208 gnd vdd FILL
XFILL_22_CLKBUF1_24 gnd vdd FILL
XFILL_74_DFFSR_219 gnd vdd FILL
XFILL_22_CLKBUF1_35 gnd vdd FILL
XFILL_18_DFFSR_30 gnd vdd FILL
XFILL_1_BUFX4_70 gnd vdd FILL
XFILL_1_BUFX4_81 gnd vdd FILL
XFILL_28_NOR3X1_18 gnd vdd FILL
XFILL_18_DFFSR_41 gnd vdd FILL
XFILL_5_CLKBUF1_17 gnd vdd FILL
XFILL_5_CLKBUF1_28 gnd vdd FILL
XFILL_1_BUFX4_92 gnd vdd FILL
XFILL_18_DFFSR_52 gnd vdd FILL
XFILL_28_NOR3X1_29 gnd vdd FILL
XFILL_18_DFFSR_63 gnd vdd FILL
XFILL_18_DFFSR_74 gnd vdd FILL
XFILL_5_CLKBUF1_39 gnd vdd FILL
XFILL_78_DFFSR_207 gnd vdd FILL
XFILL_0_AOI21X1_14 gnd vdd FILL
XFILL_18_DFFSR_85 gnd vdd FILL
XFILL_0_AOI21X1_25 gnd vdd FILL
XFILL_78_DFFSR_218 gnd vdd FILL
XFILL_13_DFFSR_140 gnd vdd FILL
XFILL_18_DFFSR_96 gnd vdd FILL
XFILL_78_DFFSR_229 gnd vdd FILL
XFILL_13_DFFSR_151 gnd vdd FILL
XFILL_0_AOI21X1_36 gnd vdd FILL
XFILL_13_DFFSR_162 gnd vdd FILL
XFILL_0_AOI21X1_47 gnd vdd FILL
XFILL_58_DFFSR_40 gnd vdd FILL
XFILL_29_NOR3X1_4 gnd vdd FILL
XFILL_0_AOI21X1_58 gnd vdd FILL
XFILL_0_AOI21X1_69 gnd vdd FILL
XFILL_13_DFFSR_173 gnd vdd FILL
XFILL_10_OAI22X1_16 gnd vdd FILL
XFILL_2_CLKBUF1_5 gnd vdd FILL
XFILL_13_DFFSR_184 gnd vdd FILL
XFILL_58_DFFSR_51 gnd vdd FILL
XFILL_10_OAI22X1_27 gnd vdd FILL
XFILL_58_DFFSR_62 gnd vdd FILL
XFILL_10_OAI22X1_38 gnd vdd FILL
XFILL_13_DFFSR_195 gnd vdd FILL
XFILL_3_NOR2X1_102 gnd vdd FILL
XFILL_58_DFFSR_73 gnd vdd FILL
XFILL_10_OAI22X1_49 gnd vdd FILL
XFILL_3_NOR2X1_113 gnd vdd FILL
XFILL_58_DFFSR_84 gnd vdd FILL
XFILL_58_DFFSR_95 gnd vdd FILL
XFILL_14_OAI21X1_18 gnd vdd FILL
XFILL_4_DFFSR_1 gnd vdd FILL
XFILL_3_NOR2X1_124 gnd vdd FILL
XFILL_14_OAI21X1_29 gnd vdd FILL
XFILL_17_DFFSR_150 gnd vdd FILL
XFILL_3_NOR2X1_135 gnd vdd FILL
XFILL_17_DFFSR_161 gnd vdd FILL
XFILL_3_NOR2X1_146 gnd vdd FILL
XFILL_3_NOR2X1_157 gnd vdd FILL
XFILL_3_NOR2X1_5 gnd vdd FILL
XFILL_17_DFFSR_172 gnd vdd FILL
XFILL_6_CLKBUF1_4 gnd vdd FILL
XFILL_3_NOR2X1_168 gnd vdd FILL
XFILL_58_0_2 gnd vdd FILL
XFILL_17_DFFSR_183 gnd vdd FILL
XFILL_3_NOR2X1_179 gnd vdd FILL
XFILL_17_DFFSR_194 gnd vdd FILL
XFILL_27_DFFSR_50 gnd vdd FILL
XFILL_27_DFFSR_61 gnd vdd FILL
XFILL_27_DFFSR_72 gnd vdd FILL
XFILL_27_DFFSR_83 gnd vdd FILL
XFILL_27_DFFSR_94 gnd vdd FILL
XFILL_27_4_0 gnd vdd FILL
XFILL_2_4_0 gnd vdd FILL
XFILL_13_NOR3X1_40 gnd vdd FILL
XFILL_20_MUX2X1_104 gnd vdd FILL
XFILL_2_MUX2X1_3 gnd vdd FILL
XFILL_13_NOR3X1_51 gnd vdd FILL
XFILL_20_MUX2X1_115 gnd vdd FILL
XFILL_67_DFFSR_60 gnd vdd FILL
XFILL_20_MUX2X1_126 gnd vdd FILL
XFILL_20_MUX2X1_137 gnd vdd FILL
XFILL_67_DFFSR_71 gnd vdd FILL
XFILL_67_DFFSR_82 gnd vdd FILL
XFILL_20_MUX2X1_148 gnd vdd FILL
XFILL_63_DFFSR_240 gnd vdd FILL
XFILL_67_DFFSR_93 gnd vdd FILL
XFILL_20_MUX2X1_159 gnd vdd FILL
XFILL_63_DFFSR_251 gnd vdd FILL
XFILL_63_DFFSR_262 gnd vdd FILL
XFILL_63_DFFSR_273 gnd vdd FILL
XFILL_3_MUX2X1_108 gnd vdd FILL
XFILL_3_MUX2X1_119 gnd vdd FILL
XFILL_39_DFFSR_3 gnd vdd FILL
XFILL_17_NOR3X1_50 gnd vdd FILL
XFILL_8_NOR2X1_202 gnd vdd FILL
XFILL_0_OAI22X1_11 gnd vdd FILL
XFILL_10_OR2X2_1 gnd vdd FILL
XFILL_0_OAI22X1_22 gnd vdd FILL
XFILL_0_OAI22X1_33 gnd vdd FILL
XFILL_67_DFFSR_250 gnd vdd FILL
XFILL_0_OAI22X1_44 gnd vdd FILL
XFILL_10_3_0 gnd vdd FILL
XFILL_67_DFFSR_261 gnd vdd FILL
XFILL_67_DFFSR_272 gnd vdd FILL
XFILL_36_DFFSR_70 gnd vdd FILL
XFILL_22_CLKBUF1_2 gnd vdd FILL
XFILL_4_OAI21X1_13 gnd vdd FILL
XFILL_4_OAI21X1_24 gnd vdd FILL
XFILL_36_DFFSR_81 gnd vdd FILL
XFILL_0_NOR2X1_12 gnd vdd FILL
XFILL_36_DFFSR_92 gnd vdd FILL
XFILL_41_DFFSR_208 gnd vdd FILL
XFILL_4_OAI21X1_35 gnd vdd FILL
XFILL_41_DFFSR_219 gnd vdd FILL
XFILL_4_OAI21X1_46 gnd vdd FILL
XFILL_0_NOR2X1_23 gnd vdd FILL
XFILL_3_OAI21X1_9 gnd vdd FILL
XFILL_0_NOR2X1_34 gnd vdd FILL
XFILL_0_NOR2X1_45 gnd vdd FILL
XFILL_0_NOR2X1_56 gnd vdd FILL
XAOI21X1_60 BUFX4_77/Y NOR2X1_28/B NOR2X1_28/Y gnd DFFSR_203/D vdd AOI21X1
XAOI21X1_71 DFFSR_149/Q NOR2X1_43/Y NOR2X1_62/Y gnd NAND3X1_85/B vdd AOI21X1
XFILL_0_NOR2X1_67 gnd vdd FILL
XFILL_0_NOR2X1_78 gnd vdd FILL
XFILL_26_CLKBUF1_1 gnd vdd FILL
XFILL_76_DFFSR_80 gnd vdd FILL
XFILL_0_NOR2X1_89 gnd vdd FILL
XFILL_4_NOR2X1_11 gnd vdd FILL
XFILL_45_DFFSR_207 gnd vdd FILL
XFILL_76_DFFSR_91 gnd vdd FILL
XFILL_4_NOR2X1_22 gnd vdd FILL
XFILL_23_DFFSR_9 gnd vdd FILL
XFILL_45_DFFSR_218 gnd vdd FILL
XFILL_7_OAI21X1_8 gnd vdd FILL
XFILL_4_NOR2X1_33 gnd vdd FILL
XFILL_45_DFFSR_229 gnd vdd FILL
XFILL_4_NOR2X1_44 gnd vdd FILL
XFILL_4_NOR2X1_55 gnd vdd FILL
XFILL_4_NOR2X1_66 gnd vdd FILL
XFILL_4_NOR2X1_77 gnd vdd FILL
XFILL_4_NOR2X1_88 gnd vdd FILL
XFILL_72_DFFSR_107 gnd vdd FILL
XFILL_11_CLKBUF1_20 gnd vdd FILL
XFILL_4_NOR2X1_99 gnd vdd FILL
XFILL_8_NOR2X1_10 gnd vdd FILL
XFILL_49_DFFSR_206 gnd vdd FILL
XFILL_8_NOR2X1_21 gnd vdd FILL
XFILL_49_DFFSR_217 gnd vdd FILL
XFILL_11_CLKBUF1_31 gnd vdd FILL
XFILL_72_DFFSR_118 gnd vdd FILL
XFILL_11_CLKBUF1_42 gnd vdd FILL
XFILL_49_DFFSR_228 gnd vdd FILL
XFILL_72_DFFSR_129 gnd vdd FILL
XFILL_8_NOR2X1_32 gnd vdd FILL
XFILL_49_0_2 gnd vdd FILL
XFILL_8_NOR2X1_43 gnd vdd FILL
XFILL_49_DFFSR_239 gnd vdd FILL
XFILL_45_DFFSR_90 gnd vdd FILL
XFILL_8_NOR2X1_54 gnd vdd FILL
XFILL_12_OAI22X1_5 gnd vdd FILL
XFILL_8_NOR2X1_65 gnd vdd FILL
XFILL_8_NOR2X1_76 gnd vdd FILL
XFILL_8_NOR2X1_87 gnd vdd FILL
XFILL_76_DFFSR_106 gnd vdd FILL
XFILL_8_NOR2X1_98 gnd vdd FILL
XFILL_76_DFFSR_117 gnd vdd FILL
XFILL_18_4_0 gnd vdd FILL
XFILL_76_DFFSR_128 gnd vdd FILL
XFILL_76_DFFSR_139 gnd vdd FILL
XFILL_16_OAI22X1_4 gnd vdd FILL
XFILL_61_7_1 gnd vdd FILL
XFILL_60_2_0 gnd vdd FILL
XFILL_26_5 gnd vdd FILL
XFILL_30_DFFSR_240 gnd vdd FILL
XFILL_30_DFFSR_251 gnd vdd FILL
XFILL_30_DFFSR_262 gnd vdd FILL
XFILL_19_4 gnd vdd FILL
XFILL_30_DFFSR_273 gnd vdd FILL
XFILL_34_DFFSR_250 gnd vdd FILL
XFILL_34_DFFSR_261 gnd vdd FILL
XFILL_34_DFFSR_272 gnd vdd FILL
XFILL_0_MUX2X1_30 gnd vdd FILL
XFILL_0_MUX2X1_41 gnd vdd FILL
XFILL_0_MUX2X1_52 gnd vdd FILL
XFILL_0_MUX2X1_63 gnd vdd FILL
XFILL_61_DFFSR_150 gnd vdd FILL
XFILL_0_MUX2X1_74 gnd vdd FILL
XFILL_61_DFFSR_161 gnd vdd FILL
XFILL_0_MUX2X1_85 gnd vdd FILL
XFILL_0_MUX2X1_96 gnd vdd FILL
XFILL_38_DFFSR_260 gnd vdd FILL
XFILL_38_DFFSR_271 gnd vdd FILL
XFILL_61_DFFSR_172 gnd vdd FILL
XFILL_61_DFFSR_183 gnd vdd FILL
XFILL_61_DFFSR_194 gnd vdd FILL
XFILL_8_NAND2X1_9 gnd vdd FILL
XFILL_12_DFFSR_207 gnd vdd FILL
XFILL_4_MUX2X1_40 gnd vdd FILL
XFILL_4_MUX2X1_51 gnd vdd FILL
XFILL_12_DFFSR_218 gnd vdd FILL
XFILL_4_MUX2X1_62 gnd vdd FILL
XFILL_4_MUX2X1_73 gnd vdd FILL
XFILL_12_DFFSR_229 gnd vdd FILL
XFILL_65_DFFSR_160 gnd vdd FILL
XFILL_4_MUX2X1_84 gnd vdd FILL
XFILL_4_MUX2X1_95 gnd vdd FILL
XFILL_65_DFFSR_171 gnd vdd FILL
XFILL_65_DFFSR_182 gnd vdd FILL
XFILL_65_DFFSR_193 gnd vdd FILL
XFILL_16_DFFSR_206 gnd vdd FILL
XFILL_10_BUFX4_16 gnd vdd FILL
XFILL_10_BUFX4_27 gnd vdd FILL
XFILL_16_DFFSR_217 gnd vdd FILL
XFILL_13_NAND3X1_6 gnd vdd FILL
XFILL_8_MUX2X1_50 gnd vdd FILL
XFILL_16_DFFSR_228 gnd vdd FILL
XFILL_8_MUX2X1_61 gnd vdd FILL
XFILL_10_BUFX4_38 gnd vdd FILL
XFILL_10_BUFX4_49 gnd vdd FILL
XFILL_8_MUX2X1_72 gnd vdd FILL
XFILL_8_MUX2X1_83 gnd vdd FILL
XFILL_16_DFFSR_239 gnd vdd FILL
XFILL_69_DFFSR_170 gnd vdd FILL
XFILL_8_MUX2X1_94 gnd vdd FILL
XFILL_69_DFFSR_181 gnd vdd FILL
XFILL_43_DFFSR_106 gnd vdd FILL
XFILL_69_DFFSR_192 gnd vdd FILL
XFILL_43_DFFSR_117 gnd vdd FILL
XFILL_43_DFFSR_128 gnd vdd FILL
XFILL_43_DFFSR_139 gnd vdd FILL
XFILL_52_7_1 gnd vdd FILL
XFILL_51_2_0 gnd vdd FILL
XFILL_47_DFFSR_105 gnd vdd FILL
XFILL_47_DFFSR_116 gnd vdd FILL
XFILL_40_DFFSR_3 gnd vdd FILL
XFILL_47_DFFSR_127 gnd vdd FILL
XFILL_8_DFFSR_2 gnd vdd FILL
XFILL_47_DFFSR_138 gnd vdd FILL
XFILL_47_DFFSR_149 gnd vdd FILL
XFILL_12_NAND3X1_14 gnd vdd FILL
XFILL_20_MUX2X1_60 gnd vdd FILL
XFILL_12_NAND3X1_25 gnd vdd FILL
XFILL_20_MUX2X1_71 gnd vdd FILL
XFILL_78_DFFSR_1 gnd vdd FILL
XFILL_12_NAND3X1_36 gnd vdd FILL
XFILL_20_MUX2X1_82 gnd vdd FILL
XFILL_20_MUX2X1_93 gnd vdd FILL
XFILL_4_INVX1_17 gnd vdd FILL
XFILL_12_NAND3X1_47 gnd vdd FILL
XFILL_12_NAND3X1_58 gnd vdd FILL
XFILL_4_INVX1_28 gnd vdd FILL
XFILL_12_NAND3X1_69 gnd vdd FILL
XFILL_32_CLKBUF1_14 gnd vdd FILL
XFILL_4_INVX1_39 gnd vdd FILL
XFILL_32_CLKBUF1_25 gnd vdd FILL
XFILL_32_CLKBUF1_36 gnd vdd FILL
XFILL_3_BUFX2_8 gnd vdd FILL
XFILL_2_BUFX4_15 gnd vdd FILL
XFILL_2_BUFX4_26 gnd vdd FILL
XFILL_62_DFFSR_7 gnd vdd FILL
XFILL_2_BUFX4_37 gnd vdd FILL
XFILL_19_DFFSR_19 gnd vdd FILL
XFILL_2_BUFX4_48 gnd vdd FILL
XFILL_2_BUFX4_59 gnd vdd FILL
XFILL_59_3_0 gnd vdd FILL
XFILL_6_0_2 gnd vdd FILL
XFILL_32_DFFSR_160 gnd vdd FILL
XFILL_32_DFFSR_171 gnd vdd FILL
XFILL_32_DFFSR_182 gnd vdd FILL
XFILL_32_DFFSR_193 gnd vdd FILL
XFILL_59_DFFSR_18 gnd vdd FILL
XFILL_59_DFFSR_29 gnd vdd FILL
XFILL_2_NAND3X1_20 gnd vdd FILL
XFILL_2_NAND3X1_31 gnd vdd FILL
XFILL_2_NAND3X1_42 gnd vdd FILL
XFILL_2_NAND3X1_53 gnd vdd FILL
XFILL_36_DFFSR_170 gnd vdd FILL
XFILL_6_NAND2X1_11 gnd vdd FILL
XFILL_2_NAND3X1_64 gnd vdd FILL
XFILL_6_NAND2X1_22 gnd vdd FILL
XFILL_2_NAND3X1_75 gnd vdd FILL
XFILL_36_DFFSR_181 gnd vdd FILL
XFILL_6_NAND2X1_33 gnd vdd FILL
XFILL_10_DFFSR_106 gnd vdd FILL
XFILL_2_BUFX4_2 gnd vdd FILL
XFILL_2_NAND3X1_86 gnd vdd FILL
XFILL_36_DFFSR_192 gnd vdd FILL
XFILL_43_7_1 gnd vdd FILL
XFILL_6_NAND2X1_44 gnd vdd FILL
XFILL_2_NAND3X1_97 gnd vdd FILL
XFILL_6_NAND2X1_55 gnd vdd FILL
XFILL_10_DFFSR_117 gnd vdd FILL
XFILL_6_NAND2X1_66 gnd vdd FILL
XFILL_42_2_0 gnd vdd FILL
XFILL_10_DFFSR_128 gnd vdd FILL
XFILL_6_NAND2X1_77 gnd vdd FILL
XFILL_10_DFFSR_139 gnd vdd FILL
XFILL_28_DFFSR_17 gnd vdd FILL
XMUX2X1_4 MUX2X1_4/A MUX2X1_4/B MUX2X1_7/S gnd MUX2X1_4/Y vdd MUX2X1
XFILL_6_NAND2X1_88 gnd vdd FILL
XFILL_28_DFFSR_28 gnd vdd FILL
XFILL_28_DFFSR_39 gnd vdd FILL
XFILL_14_DFFSR_105 gnd vdd FILL
XFILL_14_CLKBUF1_19 gnd vdd FILL
XFILL_14_DFFSR_116 gnd vdd FILL
XFILL_14_DFFSR_127 gnd vdd FILL
XFILL_14_DFFSR_138 gnd vdd FILL
XFILL_14_DFFSR_149 gnd vdd FILL
XFILL_68_DFFSR_16 gnd vdd FILL
XFILL_68_DFFSR_27 gnd vdd FILL
XFILL_68_DFFSR_38 gnd vdd FILL
XFILL_68_DFFSR_49 gnd vdd FILL
XFILL_82_DFFSR_260 gnd vdd FILL
XFILL_18_DFFSR_104 gnd vdd FILL
XFILL_82_DFFSR_271 gnd vdd FILL
XFILL_18_DFFSR_115 gnd vdd FILL
XFILL_1_INVX1_6 gnd vdd FILL
XFILL_18_DFFSR_126 gnd vdd FILL
XFILL_18_DFFSR_137 gnd vdd FILL
XFILL_18_DFFSR_148 gnd vdd FILL
XFILL_18_DFFSR_159 gnd vdd FILL
XCLKBUF1_5 BUFX4_9/Y gnd CLKBUF1_5/Y vdd CLKBUF1
XFILL_10_NOR3X1_17 gnd vdd FILL
XFILL_86_DFFSR_270 gnd vdd FILL
XFILL_10_NOR3X1_28 gnd vdd FILL
XFILL_37_DFFSR_15 gnd vdd FILL
XFILL_37_DFFSR_26 gnd vdd FILL
XFILL_37_DFFSR_37 gnd vdd FILL
XFILL_10_NOR3X1_39 gnd vdd FILL
XFILL_60_DFFSR_206 gnd vdd FILL
XFILL_37_DFFSR_48 gnd vdd FILL
XFILL_60_DFFSR_217 gnd vdd FILL
XFILL_37_DFFSR_59 gnd vdd FILL
XFILL_60_DFFSR_228 gnd vdd FILL
XFILL_60_DFFSR_239 gnd vdd FILL
XFILL_14_NOR3X1_16 gnd vdd FILL
XFILL_77_DFFSR_14 gnd vdd FILL
XFILL_14_NOR3X1_27 gnd vdd FILL
XFILL_14_NOR3X1_38 gnd vdd FILL
XFILL_77_DFFSR_25 gnd vdd FILL
XFILL_21_CLKBUF1_10 gnd vdd FILL
XFILL_21_CLKBUF1_21 gnd vdd FILL
XFILL_77_DFFSR_36 gnd vdd FILL
XFILL_14_NOR3X1_49 gnd vdd FILL
XFILL_64_DFFSR_205 gnd vdd FILL
XFILL_77_DFFSR_47 gnd vdd FILL
XFILL_21_CLKBUF1_32 gnd vdd FILL
XFILL_77_DFFSR_58 gnd vdd FILL
XFILL_64_DFFSR_216 gnd vdd FILL
XFILL_64_DFFSR_227 gnd vdd FILL
XFILL_77_DFFSR_69 gnd vdd FILL
XFILL_64_DFFSR_238 gnd vdd FILL
XFILL_0_INVX1_10 gnd vdd FILL
XFILL_0_INVX1_21 gnd vdd FILL
XFILL_64_DFFSR_249 gnd vdd FILL
XFILL_0_INVX1_32 gnd vdd FILL
XFILL_18_NOR3X1_15 gnd vdd FILL
XFILL_4_CLKBUF1_14 gnd vdd FILL
XFILL_4_CLKBUF1_25 gnd vdd FILL
XFILL_18_NOR3X1_26 gnd vdd FILL
XFILL_0_INVX1_43 gnd vdd FILL
XFILL_4_CLKBUF1_36 gnd vdd FILL
XFILL_0_INVX1_54 gnd vdd FILL
XFILL_1_AND2X2_2 gnd vdd FILL
XFILL_18_NOR3X1_37 gnd vdd FILL
XNOR2X1_203 NOR2X1_25/A NOR2X1_7/B gnd MUX2X1_22/S vdd NOR2X1
XFILL_18_NOR3X1_48 gnd vdd FILL
XFILL_0_INVX1_65 gnd vdd FILL
XFILL_68_DFFSR_204 gnd vdd FILL
XFILL_46_DFFSR_13 gnd vdd FILL
XFILL_68_DFFSR_215 gnd vdd FILL
XFILL_0_INVX1_76 gnd vdd FILL
XFILL_46_DFFSR_24 gnd vdd FILL
XFILL_68_DFFSR_226 gnd vdd FILL
XFILL_0_INVX1_87 gnd vdd FILL
XFILL_0_INVX1_98 gnd vdd FILL
XFILL_68_DFFSR_237 gnd vdd FILL
XFILL_46_DFFSR_35 gnd vdd FILL
XFILL_34_7_1 gnd vdd FILL
XFILL_31_3 gnd vdd FILL
XFILL_46_DFFSR_46 gnd vdd FILL
XFILL_68_DFFSR_248 gnd vdd FILL
XFILL_46_DFFSR_57 gnd vdd FILL
XFILL_68_DFFSR_259 gnd vdd FILL
XFILL_46_DFFSR_68 gnd vdd FILL
XFILL_33_2_0 gnd vdd FILL
XFILL_46_DFFSR_79 gnd vdd FILL
XFILL_24_2 gnd vdd FILL
XFILL_2_NOR2X1_110 gnd vdd FILL
XFILL_13_OAI21X1_15 gnd vdd FILL
XFILL_86_DFFSR_12 gnd vdd FILL
XFILL_2_NOR2X1_121 gnd vdd FILL
XFILL_13_OAI21X1_26 gnd vdd FILL
XFILL_86_DFFSR_23 gnd vdd FILL
XFILL_2_NOR2X1_132 gnd vdd FILL
XFILL_13_OAI21X1_37 gnd vdd FILL
XFILL_86_DFFSR_34 gnd vdd FILL
XFILL_17_1 gnd vdd FILL
XFILL_2_NOR2X1_143 gnd vdd FILL
XFILL_13_OAI21X1_48 gnd vdd FILL
XFILL_2_NOR2X1_154 gnd vdd FILL
XFILL_86_DFFSR_45 gnd vdd FILL
XFILL_86_DFFSR_56 gnd vdd FILL
XFILL_15_DFFSR_12 gnd vdd FILL
XFILL_2_NOR2X1_165 gnd vdd FILL
XFILL_2_NOR2X1_176 gnd vdd FILL
XFILL_86_DFFSR_67 gnd vdd FILL
XFILL_15_DFFSR_23 gnd vdd FILL
XFILL_86_DFFSR_78 gnd vdd FILL
XFILL_15_DFFSR_34 gnd vdd FILL
XFILL_86_DFFSR_89 gnd vdd FILL
XFILL_2_NOR2X1_187 gnd vdd FILL
XFILL_2_NOR2X1_198 gnd vdd FILL
XFILL_15_DFFSR_45 gnd vdd FILL
XFILL_15_DFFSR_56 gnd vdd FILL
XFILL_26_12 gnd vdd FILL
XFILL_15_DFFSR_67 gnd vdd FILL
XFILL_15_DFFSR_78 gnd vdd FILL
XFILL_15_DFFSR_89 gnd vdd FILL
XFILL_55_DFFSR_11 gnd vdd FILL
XFILL_55_DFFSR_22 gnd vdd FILL
XFILL_55_DFFSR_33 gnd vdd FILL
XFILL_26_NOR3X1_8 gnd vdd FILL
XFILL_55_DFFSR_44 gnd vdd FILL
XFILL_9_NOR2X1_19 gnd vdd FILL
XFILL_55_DFFSR_55 gnd vdd FILL
XFILL_55_DFFSR_66 gnd vdd FILL
XFILL_55_DFFSR_77 gnd vdd FILL
XFILL_55_DFFSR_88 gnd vdd FILL
XFILL_55_DFFSR_99 gnd vdd FILL
XFILL_53_DFFSR_270 gnd vdd FILL
XFILL_2_MUX2X1_105 gnd vdd FILL
XFILL_0_NOR2X1_9 gnd vdd FILL
XFILL_2_MUX2X1_116 gnd vdd FILL
XFILL_44_DFFSR_4 gnd vdd FILL
XFILL_2_MUX2X1_127 gnd vdd FILL
XFILL_2_MUX2X1_138 gnd vdd FILL
XFILL_24_DFFSR_10 gnd vdd FILL
XFILL_24_DFFSR_21 gnd vdd FILL
XFILL_2_MUX2X1_149 gnd vdd FILL
XFILL_24_DFFSR_32 gnd vdd FILL
XFILL_24_DFFSR_43 gnd vdd FILL
XFILL_24_DFFSR_54 gnd vdd FILL
XFILL_80_DFFSR_170 gnd vdd FILL
XFILL_24_DFFSR_65 gnd vdd FILL
XFILL_24_DFFSR_76 gnd vdd FILL
XFILL_3_OAI21X1_10 gnd vdd FILL
XFILL_24_DFFSR_87 gnd vdd FILL
XFILL_80_DFFSR_181 gnd vdd FILL
XFILL_24_DFFSR_98 gnd vdd FILL
XFILL_3_OAI21X1_21 gnd vdd FILL
XFILL_80_DFFSR_192 gnd vdd FILL
XFILL_31_DFFSR_205 gnd vdd FILL
XFILL_9_NOR3X1_9 gnd vdd FILL
XFILL_3_OAI21X1_32 gnd vdd FILL
XFILL_31_DFFSR_216 gnd vdd FILL
XFILL_64_DFFSR_20 gnd vdd FILL
XFILL_3_OAI21X1_43 gnd vdd FILL
XFILL_31_DFFSR_227 gnd vdd FILL
XFILL_64_DFFSR_31 gnd vdd FILL
XFILL_7_BUFX2_9 gnd vdd FILL
XFILL_64_DFFSR_42 gnd vdd FILL
XFILL_0_DFFSR_240 gnd vdd FILL
XFILL_0_DFFSR_251 gnd vdd FILL
XFILL_31_DFFSR_238 gnd vdd FILL
XFILL_64_DFFSR_53 gnd vdd FILL
XFILL_31_DFFSR_249 gnd vdd FILL
XFILL_0_DFFSR_262 gnd vdd FILL
XFILL_64_DFFSR_64 gnd vdd FILL
XFILL_0_DFFSR_273 gnd vdd FILL
XFILL_64_DFFSR_75 gnd vdd FILL
XFILL_84_DFFSR_180 gnd vdd FILL
XFILL_64_DFFSR_86 gnd vdd FILL
XFILL_84_DFFSR_191 gnd vdd FILL
XFILL_25_7_1 gnd vdd FILL
XFILL_64_DFFSR_97 gnd vdd FILL
XFILL_0_7_1 gnd vdd FILL
XFILL_35_DFFSR_204 gnd vdd FILL
XFILL_35_DFFSR_215 gnd vdd FILL
XFILL_7_DFFSR_11 gnd vdd FILL
XFILL_35_DFFSR_226 gnd vdd FILL
XFILL_24_2_0 gnd vdd FILL
XFILL_35_DFFSR_237 gnd vdd FILL
XFILL_7_DFFSR_22 gnd vdd FILL
XFILL_7_DFFSR_33 gnd vdd FILL
XFILL_4_DFFSR_250 gnd vdd FILL
XFILL_35_DFFSR_248 gnd vdd FILL
XFILL_4_DFFSR_261 gnd vdd FILL
XFILL_7_DFFSR_44 gnd vdd FILL
XFILL_7_DFFSR_55 gnd vdd FILL
XFILL_66_DFFSR_8 gnd vdd FILL
XFILL_4_DFFSR_272 gnd vdd FILL
XFILL_35_DFFSR_259 gnd vdd FILL
XFILL_33_DFFSR_30 gnd vdd FILL
XFILL_1_MUX2X1_17 gnd vdd FILL
XFILL_7_DFFSR_66 gnd vdd FILL
XFILL_33_DFFSR_41 gnd vdd FILL
XFILL_62_DFFSR_104 gnd vdd FILL
XFILL_7_DFFSR_77 gnd vdd FILL
XFILL_33_DFFSR_52 gnd vdd FILL
XFILL_1_MUX2X1_28 gnd vdd FILL
XFILL_33_DFFSR_63 gnd vdd FILL
XFILL_1_MUX2X1_39 gnd vdd FILL
XFILL_39_DFFSR_203 gnd vdd FILL
XFILL_62_DFFSR_115 gnd vdd FILL
XFILL_7_DFFSR_88 gnd vdd FILL
XFILL_7_DFFSR_99 gnd vdd FILL
XFILL_33_DFFSR_74 gnd vdd FILL
XFILL_39_DFFSR_214 gnd vdd FILL
XFILL_62_DFFSR_126 gnd vdd FILL
XFILL_39_DFFSR_225 gnd vdd FILL
XFILL_62_DFFSR_137 gnd vdd FILL
XFILL_33_DFFSR_85 gnd vdd FILL
XFILL_39_DFFSR_236 gnd vdd FILL
XFILL_62_DFFSR_148 gnd vdd FILL
XFILL_33_DFFSR_96 gnd vdd FILL
XFILL_39_DFFSR_247 gnd vdd FILL
XFILL_8_DFFSR_260 gnd vdd FILL
XFILL_62_DFFSR_159 gnd vdd FILL
XFILL_8_DFFSR_271 gnd vdd FILL
XFILL_39_DFFSR_258 gnd vdd FILL
XFILL_39_DFFSR_269 gnd vdd FILL
XFILL_5_MUX2X1_16 gnd vdd FILL
XFILL_73_DFFSR_40 gnd vdd FILL
XFILL_73_DFFSR_51 gnd vdd FILL
XFILL_66_DFFSR_103 gnd vdd FILL
XFILL_5_MUX2X1_27 gnd vdd FILL
XFILL_66_DFFSR_114 gnd vdd FILL
XFILL_73_DFFSR_62 gnd vdd FILL
XFILL_5_MUX2X1_38 gnd vdd FILL
XFILL_73_DFFSR_73 gnd vdd FILL
XFILL_5_MUX2X1_49 gnd vdd FILL
XFILL_73_DFFSR_84 gnd vdd FILL
XFILL_5_NAND3X1_19 gnd vdd FILL
XFILL_66_DFFSR_125 gnd vdd FILL
XFILL_66_DFFSR_136 gnd vdd FILL
XFILL_73_DFFSR_95 gnd vdd FILL
XFILL_66_DFFSR_147 gnd vdd FILL
XFILL_66_DFFSR_158 gnd vdd FILL
XFILL_66_DFFSR_169 gnd vdd FILL
XFILL_9_MUX2X1_15 gnd vdd FILL
XFILL_6_BUFX4_3 gnd vdd FILL
XFILL_9_MUX2X1_26 gnd vdd FILL
XFILL_9_MUX2X1_37 gnd vdd FILL
XFILL_9_MUX2X1_48 gnd vdd FILL
XFILL_13_NOR3X1_3 gnd vdd FILL
XFILL_9_MUX2X1_59 gnd vdd FILL
XFILL_13_OAI21X1_3 gnd vdd FILL
XFILL_42_DFFSR_50 gnd vdd FILL
XFILL_19_MUX2X1_130 gnd vdd FILL
XFILL_42_DFFSR_61 gnd vdd FILL
XFILL_19_MUX2X1_141 gnd vdd FILL
XFILL_10_NOR2X1_50 gnd vdd FILL
XFILL_42_DFFSR_72 gnd vdd FILL
XFILL_42_DFFSR_83 gnd vdd FILL
XFILL_10_NOR2X1_61 gnd vdd FILL
XFILL_19_MUX2X1_152 gnd vdd FILL
XFILL_19_MUX2X1_163 gnd vdd FILL
XFILL_20_DFFSR_270 gnd vdd FILL
XFILL_42_DFFSR_94 gnd vdd FILL
XFILL_10_NOR2X1_72 gnd vdd FILL
XFILL_7_3_0 gnd vdd FILL
XFILL_19_MUX2X1_174 gnd vdd FILL
XFILL_1_INVX1_210 gnd vdd FILL
XBUFX4_16 BUFX4_44/A gnd DFFSR_56/R vdd BUFX4
XFILL_10_NOR2X1_83 gnd vdd FILL
XBUFX4_27 BUFX4_47/A gnd DFFSR_58/R vdd BUFX4
XFILL_19_MUX2X1_185 gnd vdd FILL
XFILL_10_NOR2X1_94 gnd vdd FILL
XFILL_1_INVX1_221 gnd vdd FILL
XBUFX4_38 BUFX4_47/A gnd DFFSR_23/R vdd BUFX4
XBUFX4_49 BUFX4_62/Y gnd DFFSR_98/R vdd BUFX4
XFILL_82_DFFSR_60 gnd vdd FILL
XFILL_82_DFFSR_71 gnd vdd FILL
XFILL_82_DFFSR_82 gnd vdd FILL
XFILL_82_DFFSR_93 gnd vdd FILL
XFILL_11_DFFSR_60 gnd vdd FILL
XFILL_21_MUX2X1_14 gnd vdd FILL
XFILL_5_INVX1_220 gnd vdd FILL
XFILL_21_MUX2X1_25 gnd vdd FILL
XFILL_11_DFFSR_71 gnd vdd FILL
XFILL_5_INVX1_7 gnd vdd FILL
XFILL_11_DFFSR_82 gnd vdd FILL
XFILL_21_MUX2X1_36 gnd vdd FILL
XFILL_11_DFFSR_93 gnd vdd FILL
XFILL_21_MUX2X1_47 gnd vdd FILL
XFILL_21_MUX2X1_58 gnd vdd FILL
XFILL_21_MUX2X1_69 gnd vdd FILL
XFILL_16_7_1 gnd vdd FILL
XFILL_22_NOR3X1_1 gnd vdd FILL
XFILL_15_2_0 gnd vdd FILL
XFILL_51_DFFSR_180 gnd vdd FILL
XFILL_51_DFFSR_191 gnd vdd FILL
XFILL_51_DFFSR_70 gnd vdd FILL
XFILL_51_DFFSR_81 gnd vdd FILL
XFILL_51_DFFSR_92 gnd vdd FILL
XFILL_55_DFFSR_190 gnd vdd FILL
XFILL_20_DFFSR_80 gnd vdd FILL
XFILL_20_DFFSR_91 gnd vdd FILL
XFILL_9_MUX2X1_180 gnd vdd FILL
XFILL_9_INVX8_1 gnd vdd FILL
XFILL_5_NOR3X1_2 gnd vdd FILL
XFILL_9_MUX2X1_191 gnd vdd FILL
XFILL_33_DFFSR_103 gnd vdd FILL
XFILL_33_DFFSR_114 gnd vdd FILL
XFILL_10_NAND2X1_5 gnd vdd FILL
XFILL_33_DFFSR_125 gnd vdd FILL
XFILL_33_DFFSR_136 gnd vdd FILL
XFILL_2_DFFSR_160 gnd vdd FILL
XFILL_33_DFFSR_147 gnd vdd FILL
XFILL_33_DFFSR_158 gnd vdd FILL
XFILL_2_DFFSR_171 gnd vdd FILL
XFILL_33_DFFSR_169 gnd vdd FILL
XFILL_60_DFFSR_90 gnd vdd FILL
XFILL_2_DFFSR_182 gnd vdd FILL
XFILL_2_DFFSR_193 gnd vdd FILL
XFILL_37_DFFSR_102 gnd vdd FILL
XFILL_37_DFFSR_113 gnd vdd FILL
XFILL_37_DFFSR_124 gnd vdd FILL
XFILL_5_NOR2X1_109 gnd vdd FILL
XFILL_37_DFFSR_135 gnd vdd FILL
XFILL_26_DFFSR_1 gnd vdd FILL
XFILL_37_DFFSR_146 gnd vdd FILL
XFILL_11_NAND3X1_11 gnd vdd FILL
XFILL_37_DFFSR_157 gnd vdd FILL
XFILL_6_DFFSR_170 gnd vdd FILL
XFILL_11_NAND3X1_22 gnd vdd FILL
XFILL_83_DFFSR_2 gnd vdd FILL
XFILL_37_DFFSR_168 gnd vdd FILL
XFILL_3_DFFSR_70 gnd vdd FILL
XFILL_11_NAND3X1_33 gnd vdd FILL
XFILL_6_DFFSR_181 gnd vdd FILL
XFILL_11_NAND3X1_44 gnd vdd FILL
XFILL_37_DFFSR_179 gnd vdd FILL
XFILL_10_MUX2X1_90 gnd vdd FILL
XFILL_3_DFFSR_81 gnd vdd FILL
XFILL_6_DFFSR_192 gnd vdd FILL
XFILL_11_NAND3X1_55 gnd vdd FILL
XFILL_3_DFFSR_92 gnd vdd FILL
XFILL_31_CLKBUF1_11 gnd vdd FILL
XFILL_11_NAND3X1_66 gnd vdd FILL
XFILL_66_6_1 gnd vdd FILL
XFILL_31_CLKBUF1_22 gnd vdd FILL
XFILL_11_NAND3X1_77 gnd vdd FILL
XFILL_11_NAND3X1_88 gnd vdd FILL
XFILL_65_1_0 gnd vdd FILL
XFILL_31_CLKBUF1_33 gnd vdd FILL
XFILL_11_NAND3X1_99 gnd vdd FILL
XFILL_83_DFFSR_203 gnd vdd FILL
XFILL_83_DFFSR_214 gnd vdd FILL
XFILL_83_DFFSR_225 gnd vdd FILL
XFILL_83_DFFSR_236 gnd vdd FILL
XFILL_10_DFFSR_7 gnd vdd FILL
XFILL_83_DFFSR_247 gnd vdd FILL
XFILL_83_DFFSR_258 gnd vdd FILL
XFILL_83_DFFSR_269 gnd vdd FILL
XFILL_48_DFFSR_5 gnd vdd FILL
XFILL_87_DFFSR_202 gnd vdd FILL
XFILL_87_DFFSR_213 gnd vdd FILL
XFILL_87_DFFSR_224 gnd vdd FILL
XFILL_87_DFFSR_235 gnd vdd FILL
XFILL_14_AOI21X1_9 gnd vdd FILL
XFILL_2_OAI22X1_18 gnd vdd FILL
XFILL_2_OAI22X1_29 gnd vdd FILL
XFILL_87_DFFSR_246 gnd vdd FILL
XFILL_87_DFFSR_257 gnd vdd FILL
XFILL_87_DFFSR_268 gnd vdd FILL
XFILL_22_DFFSR_190 gnd vdd FILL
XFILL_15_AOI22X1_11 gnd vdd FILL
XFILL_3_INVX1_130 gnd vdd FILL
XFILL_3_INVX1_141 gnd vdd FILL
XFILL_3_INVX1_152 gnd vdd FILL
XFILL_3_INVX1_163 gnd vdd FILL
XFILL_1_NAND3X1_50 gnd vdd FILL
XFILL_3_INVX1_174 gnd vdd FILL
XFILL_1_NAND3X1_61 gnd vdd FILL
XFILL_3_INVX1_185 gnd vdd FILL
XFILL_1_NAND3X1_72 gnd vdd FILL
XFILL_3_INVX1_196 gnd vdd FILL
XFILL_5_NAND2X1_30 gnd vdd FILL
XFILL_5_NAND2X1_41 gnd vdd FILL
XFILL_1_NAND3X1_83 gnd vdd FILL
XFILL_1_NAND3X1_94 gnd vdd FILL
XFILL_5_NAND2X1_52 gnd vdd FILL
XFILL_5_NAND2X1_63 gnd vdd FILL
XFILL_7_INVX1_140 gnd vdd FILL
XFILL_7_INVX1_151 gnd vdd FILL
XFILL_5_NAND2X1_74 gnd vdd FILL
XFILL_7_INVX1_162 gnd vdd FILL
XFILL_5_NAND2X1_85 gnd vdd FILL
XFILL_5_NAND2X1_96 gnd vdd FILL
XFILL_7_INVX1_173 gnd vdd FILL
XFILL_7_INVX1_184 gnd vdd FILL
XFILL_7_INVX1_195 gnd vdd FILL
XFILL_13_CLKBUF1_16 gnd vdd FILL
XFILL_13_CLKBUF1_27 gnd vdd FILL
XFILL_13_CLKBUF1_38 gnd vdd FILL
XFILL_1_OAI22X1_3 gnd vdd FILL
XFILL_57_6_1 gnd vdd FILL
XFILL_56_1_0 gnd vdd FILL
XFILL_11_NOR2X1_101 gnd vdd FILL
XFILL_5_OAI22X1_2 gnd vdd FILL
XFILL_11_NOR2X1_112 gnd vdd FILL
XFILL_11_NOR2X1_123 gnd vdd FILL
XFILL_11_NOR2X1_134 gnd vdd FILL
XFILL_11_NOR2X1_145 gnd vdd FILL
XFILL_11_NOR2X1_156 gnd vdd FILL
XFILL_11_NOR2X1_167 gnd vdd FILL
XFILL_11_NOR2X1_178 gnd vdd FILL
XFILL_50_DFFSR_203 gnd vdd FILL
XFILL_11_NOR2X1_189 gnd vdd FILL
XFILL_50_DFFSR_214 gnd vdd FILL
XFILL_9_OAI22X1_1 gnd vdd FILL
XFILL_50_DFFSR_225 gnd vdd FILL
XFILL_9_AOI21X1_30 gnd vdd FILL
XFILL_9_AOI21X1_41 gnd vdd FILL
XFILL_40_5_1 gnd vdd FILL
XFILL_50_DFFSR_236 gnd vdd FILL
XFILL_50_DFFSR_247 gnd vdd FILL
XFILL_9_AOI21X1_52 gnd vdd FILL
XFILL_50_DFFSR_258 gnd vdd FILL
XFILL_19_OAI22X1_10 gnd vdd FILL
XFILL_50_DFFSR_269 gnd vdd FILL
XFILL_9_AOI21X1_63 gnd vdd FILL
XFILL_19_OAI22X1_21 gnd vdd FILL
XFILL_9_AOI21X1_74 gnd vdd FILL
XFILL_19_OAI22X1_32 gnd vdd FILL
XFILL_54_DFFSR_202 gnd vdd FILL
XFILL_19_OAI22X1_43 gnd vdd FILL
XFILL_54_DFFSR_213 gnd vdd FILL
XFILL_20_CLKBUF1_40 gnd vdd FILL
XFILL_54_DFFSR_224 gnd vdd FILL
XFILL_54_DFFSR_235 gnd vdd FILL
XFILL_54_DFFSR_246 gnd vdd FILL
XFILL_3_CLKBUF1_11 gnd vdd FILL
XFILL_54_DFFSR_257 gnd vdd FILL
XFILL_3_CLKBUF1_22 gnd vdd FILL
XFILL_54_DFFSR_268 gnd vdd FILL
XFILL_3_CLKBUF1_33 gnd vdd FILL
XFILL_81_DFFSR_102 gnd vdd FILL
XFILL_58_DFFSR_201 gnd vdd FILL
XFILL_81_DFFSR_113 gnd vdd FILL
XFILL_11_MUX2X1_107 gnd vdd FILL
XFILL_34_DFFSR_19 gnd vdd FILL
XFILL_11_MUX2X1_118 gnd vdd FILL
XFILL_58_DFFSR_212 gnd vdd FILL
XFILL_81_DFFSR_124 gnd vdd FILL
XFILL_58_DFFSR_223 gnd vdd FILL
XFILL_11_MUX2X1_129 gnd vdd FILL
XFILL_58_DFFSR_234 gnd vdd FILL
XFILL_81_DFFSR_135 gnd vdd FILL
XFILL_81_DFFSR_146 gnd vdd FILL
XFILL_58_DFFSR_245 gnd vdd FILL
XFILL_81_DFFSR_157 gnd vdd FILL
XFILL_81_DFFSR_168 gnd vdd FILL
XFILL_58_DFFSR_256 gnd vdd FILL
XFILL_58_DFFSR_267 gnd vdd FILL
XFILL_81_DFFSR_179 gnd vdd FILL
XFILL_13_CLKBUF1_8 gnd vdd FILL
XFILL_1_DFFSR_205 gnd vdd FILL
XFILL_85_DFFSR_101 gnd vdd FILL
XFILL_1_DFFSR_216 gnd vdd FILL
XFILL_74_DFFSR_18 gnd vdd FILL
XFILL_85_DFFSR_112 gnd vdd FILL
XFILL_1_DFFSR_227 gnd vdd FILL
XFILL_12_OAI21X1_12 gnd vdd FILL
XFILL_85_DFFSR_123 gnd vdd FILL
XFILL_74_DFFSR_29 gnd vdd FILL
XFILL_12_OAI21X1_23 gnd vdd FILL
XFILL_85_DFFSR_134 gnd vdd FILL
XFILL_1_DFFSR_238 gnd vdd FILL
XFILL_12_OAI21X1_34 gnd vdd FILL
XFILL_85_DFFSR_145 gnd vdd FILL
XFILL_1_DFFSR_249 gnd vdd FILL
XFILL_1_NOR2X1_140 gnd vdd FILL
XFILL_12_OAI21X1_45 gnd vdd FILL
XFILL_85_DFFSR_156 gnd vdd FILL
XFILL_17_MUX2X1_8 gnd vdd FILL
XFILL_1_NOR2X1_151 gnd vdd FILL
XFILL_1_NOR2X1_162 gnd vdd FILL
XFILL_85_DFFSR_167 gnd vdd FILL
XFILL_85_DFFSR_178 gnd vdd FILL
XFILL_1_NOR2X1_173 gnd vdd FILL
XFILL_17_CLKBUF1_7 gnd vdd FILL
XFILL_1_NOR2X1_184 gnd vdd FILL
XFILL_85_DFFSR_189 gnd vdd FILL
XFILL_5_DFFSR_204 gnd vdd FILL
XFILL_2_NAND3X1_4 gnd vdd FILL
XFILL_5_DFFSR_215 gnd vdd FILL
XFILL_48_6_1 gnd vdd FILL
XFILL_1_NOR2X1_195 gnd vdd FILL
XFILL_8_BUFX4_30 gnd vdd FILL
XFILL_5_DFFSR_226 gnd vdd FILL
XFILL_8_BUFX4_41 gnd vdd FILL
XFILL_5_DFFSR_237 gnd vdd FILL
XFILL_47_1_0 gnd vdd FILL
XFILL_8_BUFX4_52 gnd vdd FILL
XFILL_5_DFFSR_248 gnd vdd FILL
XFILL_8_BUFX4_63 gnd vdd FILL
XFILL_13_BUFX4_102 gnd vdd FILL
XFILL_43_DFFSR_17 gnd vdd FILL
XFILL_5_DFFSR_259 gnd vdd FILL
XFILL_43_DFFSR_28 gnd vdd FILL
XFILL_8_BUFX4_74 gnd vdd FILL
XFILL_8_BUFX4_85 gnd vdd FILL
XFILL_8_BUFX4_96 gnd vdd FILL
XFILL_43_DFFSR_39 gnd vdd FILL
XFILL_6_NAND3X1_3 gnd vdd FILL
XFILL_9_DFFSR_203 gnd vdd FILL
XFILL_9_DFFSR_214 gnd vdd FILL
XFILL_9_DFFSR_225 gnd vdd FILL
XFILL_9_DFFSR_236 gnd vdd FILL
XFILL_9_DFFSR_247 gnd vdd FILL
XFILL_83_DFFSR_16 gnd vdd FILL
XFILL_9_DFFSR_258 gnd vdd FILL
XFILL_9_DFFSR_269 gnd vdd FILL
XFILL_83_DFFSR_27 gnd vdd FILL
XFILL_83_DFFSR_38 gnd vdd FILL
XFILL_1_MUX2X1_102 gnd vdd FILL
XFILL_1_MUX2X1_113 gnd vdd FILL
XFILL_83_DFFSR_49 gnd vdd FILL
XFILL_1_MUX2X1_124 gnd vdd FILL
XFILL_12_DFFSR_16 gnd vdd FILL
XFILL_1_MUX2X1_135 gnd vdd FILL
XFILL_12_DFFSR_27 gnd vdd FILL
XFILL_31_5_1 gnd vdd FILL
XFILL_1_MUX2X1_146 gnd vdd FILL
XFILL_12_DFFSR_38 gnd vdd FILL
XFILL_12_DFFSR_49 gnd vdd FILL
XFILL_30_0_0 gnd vdd FILL
XFILL_1_MUX2X1_157 gnd vdd FILL
XFILL_87_DFFSR_3 gnd vdd FILL
XFILL_1_MUX2X1_168 gnd vdd FILL
XFILL_1_MUX2X1_179 gnd vdd FILL
XFILL_52_DFFSR_15 gnd vdd FILL
XFILL_21_DFFSR_202 gnd vdd FILL
XFILL_52_DFFSR_26 gnd vdd FILL
XFILL_21_DFFSR_213 gnd vdd FILL
XFILL_52_DFFSR_37 gnd vdd FILL
XFILL_11_NOR2X1_15 gnd vdd FILL
XFILL_2_OAI21X1_40 gnd vdd FILL
XFILL_52_DFFSR_48 gnd vdd FILL
XFILL_21_DFFSR_224 gnd vdd FILL
XFILL_11_NOR2X1_26 gnd vdd FILL
XFILL_21_DFFSR_235 gnd vdd FILL
XFILL_2_AOI22X1_9 gnd vdd FILL
XFILL_11_NOR2X1_37 gnd vdd FILL
XFILL_52_DFFSR_59 gnd vdd FILL
XFILL_21_DFFSR_246 gnd vdd FILL
XFILL_11_NOR2X1_48 gnd vdd FILL
XFILL_11_NOR2X1_59 gnd vdd FILL
XFILL_21_DFFSR_257 gnd vdd FILL
XFILL_21_DFFSR_268 gnd vdd FILL
XFILL_2_INVX1_208 gnd vdd FILL
XFILL_25_DFFSR_201 gnd vdd FILL
XFILL_2_INVX1_219 gnd vdd FILL
XFILL_9_MUX2X1_7 gnd vdd FILL
XFILL_25_DFFSR_212 gnd vdd FILL
XFILL_25_DFFSR_223 gnd vdd FILL
XFILL_25_DFFSR_234 gnd vdd FILL
XFILL_14_DFFSR_8 gnd vdd FILL
XFILL_6_AOI22X1_8 gnd vdd FILL
XFILL_21_DFFSR_14 gnd vdd FILL
XFILL_25_DFFSR_245 gnd vdd FILL
XFILL_71_DFFSR_9 gnd vdd FILL
XFILL_21_DFFSR_25 gnd vdd FILL
XFILL_21_DFFSR_36 gnd vdd FILL
XFILL_25_DFFSR_256 gnd vdd FILL
XFILL_25_DFFSR_267 gnd vdd FILL
XFILL_21_DFFSR_47 gnd vdd FILL
XFILL_21_DFFSR_58 gnd vdd FILL
XFILL_6_INVX1_207 gnd vdd FILL
XFILL_52_DFFSR_101 gnd vdd FILL
XFILL_29_DFFSR_200 gnd vdd FILL
XFILL_12_BUFX4_90 gnd vdd FILL
XFILL_21_DFFSR_69 gnd vdd FILL
XFILL_52_DFFSR_112 gnd vdd FILL
XFILL_6_INVX1_218 gnd vdd FILL
XFILL_29_DFFSR_211 gnd vdd FILL
XFILL_52_DFFSR_123 gnd vdd FILL
XFILL_29_DFFSR_222 gnd vdd FILL
XFILL_52_DFFSR_134 gnd vdd FILL
XFILL_61_DFFSR_13 gnd vdd FILL
XFILL_29_DFFSR_233 gnd vdd FILL
XFILL_52_DFFSR_145 gnd vdd FILL
XFILL_29_DFFSR_244 gnd vdd FILL
XFILL_52_DFFSR_156 gnd vdd FILL
XFILL_61_DFFSR_24 gnd vdd FILL
XFILL_61_DFFSR_35 gnd vdd FILL
XFILL_39_6_1 gnd vdd FILL
XFILL_29_DFFSR_255 gnd vdd FILL
XFILL_52_DFFSR_167 gnd vdd FILL
XFILL_61_DFFSR_46 gnd vdd FILL
XFILL_29_DFFSR_266 gnd vdd FILL
XFILL_52_DFFSR_178 gnd vdd FILL
XFILL_61_DFFSR_57 gnd vdd FILL
XFILL_38_1_0 gnd vdd FILL
XFILL_61_DFFSR_68 gnd vdd FILL
XFILL_56_DFFSR_100 gnd vdd FILL
XFILL_52_DFFSR_189 gnd vdd FILL
XFILL_56_DFFSR_111 gnd vdd FILL
XFILL_4_NAND3X1_16 gnd vdd FILL
XFILL_61_DFFSR_79 gnd vdd FILL
XFILL_56_DFFSR_122 gnd vdd FILL
XFILL_56_DFFSR_133 gnd vdd FILL
XFILL_4_NAND3X1_27 gnd vdd FILL
XFILL_56_DFFSR_144 gnd vdd FILL
XFILL_4_NAND3X1_38 gnd vdd FILL
XFILL_56_DFFSR_155 gnd vdd FILL
XFILL_4_NAND3X1_49 gnd vdd FILL
XFILL_56_DFFSR_166 gnd vdd FILL
XFILL_4_DFFSR_15 gnd vdd FILL
XFILL_56_DFFSR_177 gnd vdd FILL
XFILL_4_DFFSR_26 gnd vdd FILL
XFILL_8_NAND2X1_18 gnd vdd FILL
XFILL_30_DFFSR_12 gnd vdd FILL
XFILL_4_DFFSR_37 gnd vdd FILL
XFILL_8_NAND2X1_29 gnd vdd FILL
XFILL_56_DFFSR_188 gnd vdd FILL
XFILL_4_DFFSR_48 gnd vdd FILL
XFILL_30_DFFSR_23 gnd vdd FILL
XFILL_56_DFFSR_199 gnd vdd FILL
XFILL_4_DFFSR_59 gnd vdd FILL
XFILL_30_DFFSR_34 gnd vdd FILL
XFILL_30_DFFSR_45 gnd vdd FILL
XFILL_30_DFFSR_56 gnd vdd FILL
XFILL_30_DFFSR_67 gnd vdd FILL
XFILL_30_DFFSR_78 gnd vdd FILL
XFILL_22_5_1 gnd vdd FILL
XFILL_30_DFFSR_89 gnd vdd FILL
XFILL_6_INVX1_80 gnd vdd FILL
XFILL_6_INVX1_91 gnd vdd FILL
XFILL_70_DFFSR_11 gnd vdd FILL
XFILL_3_DFFSR_103 gnd vdd FILL
XFILL_18_MUX2X1_160 gnd vdd FILL
XFILL_70_DFFSR_22 gnd vdd FILL
XFILL_3_DFFSR_114 gnd vdd FILL
XFILL_18_MUX2X1_171 gnd vdd FILL
XFILL_21_0_0 gnd vdd FILL
XFILL_18_MUX2X1_182 gnd vdd FILL
XFILL_70_DFFSR_33 gnd vdd FILL
XFILL_3_DFFSR_125 gnd vdd FILL
XFILL_3_DFFSR_136 gnd vdd FILL
XFILL_13_MUX2X1_1 gnd vdd FILL
XFILL_18_MUX2X1_193 gnd vdd FILL
XFILL_70_DFFSR_44 gnd vdd FILL
XFILL_70_DFFSR_55 gnd vdd FILL
XFILL_3_DFFSR_147 gnd vdd FILL
XFILL_3_DFFSR_158 gnd vdd FILL
XFILL_70_DFFSR_66 gnd vdd FILL
XFILL_70_DFFSR_77 gnd vdd FILL
XFILL_3_DFFSR_169 gnd vdd FILL
XFILL_70_DFFSR_88 gnd vdd FILL
XFILL_7_DFFSR_102 gnd vdd FILL
XFILL_70_DFFSR_99 gnd vdd FILL
XFILL_11_MUX2X1_11 gnd vdd FILL
XFILL_7_DFFSR_113 gnd vdd FILL
XFILL_7_DFFSR_124 gnd vdd FILL
XFILL_11_MUX2X1_22 gnd vdd FILL
XFILL_7_DFFSR_135 gnd vdd FILL
XFILL_11_MUX2X1_33 gnd vdd FILL
XDFFSR_160 DFFSR_160/Q DFFSR_99/CLK DFFSR_89/R vdd DFFSR_160/D gnd vdd DFFSR
XFILL_7_DFFSR_146 gnd vdd FILL
XBUFX4_1 BUFX4_2/A gnd BUFX4_1/Y vdd BUFX4
XFILL_11_MUX2X1_44 gnd vdd FILL
XFILL_7_DFFSR_157 gnd vdd FILL
XFILL_11_MUX2X1_55 gnd vdd FILL
XDFFSR_171 INVX1_79/A CLKBUF1_34/Y BUFX4_23/Y vdd MUX2X1_24/Y gnd vdd DFFSR
XFILL_11_MUX2X1_66 gnd vdd FILL
XFILL_7_DFFSR_168 gnd vdd FILL
XDFFSR_182 INVX1_196/A DFFSR_64/CLK DFFSR_69/R vdd DFFSR_182/D gnd vdd DFFSR
XFILL_11_MUX2X1_77 gnd vdd FILL
XFILL_7_DFFSR_179 gnd vdd FILL
XDFFSR_193 DFFSR_194/D CLKBUF1_24/Y DFFSR_1/R vdd next gnd vdd DFFSR
XFILL_10_NOR3X1_7 gnd vdd FILL
XFILL_11_MUX2X1_88 gnd vdd FILL
XFILL_11_MUX2X1_99 gnd vdd FILL
XFILL_15_MUX2X1_10 gnd vdd FILL
XFILL_15_MUX2X1_21 gnd vdd FILL
XFILL_15_MUX2X1_32 gnd vdd FILL
XFILL_15_MUX2X1_43 gnd vdd FILL
XFILL_15_MUX2X1_54 gnd vdd FILL
XFILL_15_MUX2X1_65 gnd vdd FILL
XFILL_15_MUX2X1_76 gnd vdd FILL
XFILL_3_NOR3X1_14 gnd vdd FILL
XFILL_15_MUX2X1_87 gnd vdd FILL
XFILL_3_NOR3X1_25 gnd vdd FILL
XFILL_3_NOR3X1_36 gnd vdd FILL
XFILL_15_MUX2X1_98 gnd vdd FILL
XFILL_3_NOR3X1_47 gnd vdd FILL
XFILL_19_MUX2X1_20 gnd vdd FILL
XFILL_19_MUX2X1_31 gnd vdd FILL
XFILL_23_CLKBUF1_17 gnd vdd FILL
XFILL_23_CLKBUF1_28 gnd vdd FILL
XFILL_19_MUX2X1_42 gnd vdd FILL
XFILL_5_6_1 gnd vdd FILL
XFILL_19_MUX2X1_53 gnd vdd FILL
XFILL_6_NOR2X1_2 gnd vdd FILL
XFILL_23_CLKBUF1_39 gnd vdd FILL
XFILL_19_MUX2X1_64 gnd vdd FILL
XFILL_4_1_0 gnd vdd FILL
XFILL_29_1_0 gnd vdd FILL
XFILL_19_MUX2X1_75 gnd vdd FILL
XFILL_7_NOR3X1_13 gnd vdd FILL
XFILL_19_MUX2X1_86 gnd vdd FILL
XFILL_7_NOR3X1_24 gnd vdd FILL
XFILL_0_INVX1_107 gnd vdd FILL
XFILL_19_MUX2X1_97 gnd vdd FILL
XFILL_7_NOR3X1_35 gnd vdd FILL
XFILL_7_NOR3X1_46 gnd vdd FILL
XFILL_0_INVX1_118 gnd vdd FILL
XFILL_23_DFFSR_100 gnd vdd FILL
XFILL_23_DFFSR_111 gnd vdd FILL
XFILL_0_INVX1_129 gnd vdd FILL
XFILL_23_DFFSR_122 gnd vdd FILL
XFILL_1_AOI21X1_18 gnd vdd FILL
XFILL_23_DFFSR_133 gnd vdd FILL
XFILL_1_AOI21X1_29 gnd vdd FILL
XFILL_23_DFFSR_144 gnd vdd FILL
XFILL_23_DFFSR_155 gnd vdd FILL
XFILL_23_DFFSR_166 gnd vdd FILL
XFILL_23_DFFSR_177 gnd vdd FILL
XFILL_4_INVX1_106 gnd vdd FILL
XFILL_4_INVX1_117 gnd vdd FILL
XFILL_23_DFFSR_188 gnd vdd FILL
XFILL_27_DFFSR_110 gnd vdd FILL
XFILL_23_DFFSR_199 gnd vdd FILL
XFILL_4_NOR2X1_106 gnd vdd FILL
XFILL_4_INVX1_128 gnd vdd FILL
XFILL_13_5_1 gnd vdd FILL
XFILL_27_DFFSR_121 gnd vdd FILL
XFILL_27_DFFSR_132 gnd vdd FILL
XFILL_4_INVX1_139 gnd vdd FILL
XFILL_4_NOR2X1_117 gnd vdd FILL
XFILL_4_NOR2X1_128 gnd vdd FILL
XFILL_31_DFFSR_2 gnd vdd FILL
XFILL_27_DFFSR_143 gnd vdd FILL
XFILL_12_0_0 gnd vdd FILL
XFILL_27_DFFSR_154 gnd vdd FILL
XFILL_4_NOR2X1_139 gnd vdd FILL
XFILL_27_DFFSR_165 gnd vdd FILL
XFILL_10_NAND3X1_30 gnd vdd FILL
XINVX4_1 INVX4_1/A gnd INVX4_1/Y vdd INVX4
XFILL_10_NAND3X1_41 gnd vdd FILL
XFILL_27_DFFSR_176 gnd vdd FILL
XFILL_10_NAND3X1_52 gnd vdd FILL
XFILL_27_DFFSR_187 gnd vdd FILL
XFILL_27_DFFSR_198 gnd vdd FILL
XFILL_10_NAND3X1_63 gnd vdd FILL
XFILL_10_NAND3X1_74 gnd vdd FILL
XFILL_30_CLKBUF1_30 gnd vdd FILL
XFILL_10_NAND3X1_85 gnd vdd FILL
XFILL_2_NOR3X1_6 gnd vdd FILL
XFILL_10_NAND3X1_96 gnd vdd FILL
XFILL_30_CLKBUF1_41 gnd vdd FILL
XFILL_23_NOR3X1_11 gnd vdd FILL
XFILL_23_NOR3X1_22 gnd vdd FILL
XFILL_23_NOR3X1_33 gnd vdd FILL
XFILL_23_NOR3X1_44 gnd vdd FILL
XFILL_73_DFFSR_200 gnd vdd FILL
XFILL_21_MUX2X1_108 gnd vdd FILL
XFILL_21_MUX2X1_119 gnd vdd FILL
XFILL_73_DFFSR_211 gnd vdd FILL
XFILL_73_DFFSR_222 gnd vdd FILL
XFILL_73_DFFSR_233 gnd vdd FILL
XFILL_0_DFFSR_30 gnd vdd FILL
XFILL_73_DFFSR_244 gnd vdd FILL
XFILL_27_NOR3X1_10 gnd vdd FILL
XFILL_0_DFFSR_41 gnd vdd FILL
XFILL_73_DFFSR_255 gnd vdd FILL
XFILL_0_DFFSR_52 gnd vdd FILL
XFILL_0_DFFSR_63 gnd vdd FILL
XFILL_53_DFFSR_6 gnd vdd FILL
XFILL_73_DFFSR_266 gnd vdd FILL
XFILL_27_NOR3X1_21 gnd vdd FILL
XFILL_0_DFFSR_74 gnd vdd FILL
XFILL_27_NOR3X1_32 gnd vdd FILL
XFILL_7_4 gnd vdd FILL
XFILL_27_NOR3X1_43 gnd vdd FILL
XFILL_0_DFFSR_85 gnd vdd FILL
XFILL_77_DFFSR_210 gnd vdd FILL
XFILL_0_DFFSR_96 gnd vdd FILL
XFILL_9_NOR2X1_206 gnd vdd FILL
XFILL_77_DFFSR_221 gnd vdd FILL
XFILL_1_OAI22X1_15 gnd vdd FILL
XFILL_77_DFFSR_232 gnd vdd FILL
XFILL_77_DFFSR_243 gnd vdd FILL
XFILL_1_OAI22X1_26 gnd vdd FILL
XFILL_63_6 gnd vdd FILL
XFILL_77_DFFSR_254 gnd vdd FILL
XFILL_1_OAI22X1_37 gnd vdd FILL
XFILL_77_DFFSR_265 gnd vdd FILL
XFILL_1_OAI22X1_48 gnd vdd FILL
XFILL_5_OAI21X1_17 gnd vdd FILL
XFILL_32_CLKBUF1_6 gnd vdd FILL
XFILL_56_5 gnd vdd FILL
XFILL_5_OAI21X1_28 gnd vdd FILL
XFILL_5_OAI21X1_39 gnd vdd FILL
XFILL_63_4_1 gnd vdd FILL
XFILL_0_NAND3X1_80 gnd vdd FILL
XFILL_0_NAND3X1_91 gnd vdd FILL
XFILL_4_NAND2X1_60 gnd vdd FILL
XFILL_18_DFFSR_9 gnd vdd FILL
XFILL_4_NAND2X1_71 gnd vdd FILL
XFILL_4_NAND2X1_82 gnd vdd FILL
XFILL_4_NAND2X1_93 gnd vdd FILL
XFILL_9_BUFX4_19 gnd vdd FILL
XFILL_12_CLKBUF1_13 gnd vdd FILL
XFILL_12_CLKBUF1_24 gnd vdd FILL
XFILL_12_CLKBUF1_35 gnd vdd FILL
XFILL_10_NOR2X1_120 gnd vdd FILL
XFILL_10_NOR2X1_131 gnd vdd FILL
XFILL_10_NOR2X1_142 gnd vdd FILL
XFILL_10_NOR2X1_153 gnd vdd FILL
XFILL_10_NOR2X1_164 gnd vdd FILL
XFILL_40_DFFSR_200 gnd vdd FILL
XFILL_10_NOR2X1_175 gnd vdd FILL
XFILL_40_DFFSR_211 gnd vdd FILL
XFILL_10_NOR2X1_186 gnd vdd FILL
XFILL_40_DFFSR_222 gnd vdd FILL
XFILL_10_NOR2X1_197 gnd vdd FILL
XFILL_2_OAI21X1_1 gnd vdd FILL
XFILL_40_DFFSR_233 gnd vdd FILL
XFILL_40_DFFSR_244 gnd vdd FILL
XFILL_40_DFFSR_255 gnd vdd FILL
XFILL_8_AOI21X1_60 gnd vdd FILL
XFILL_40_DFFSR_266 gnd vdd FILL
XNAND3X1_4 NOR2X1_91/Y NOR3X1_35/Y NOR2X1_84/Y gnd NAND3X1_4/Y vdd NAND3X1
XFILL_8_AOI21X1_71 gnd vdd FILL
XFILL_18_OAI22X1_40 gnd vdd FILL
XFILL_18_OAI22X1_51 gnd vdd FILL
XFILL_44_DFFSR_210 gnd vdd FILL
XFILL_44_DFFSR_221 gnd vdd FILL
XFILL_44_DFFSR_232 gnd vdd FILL
XFILL_44_DFFSR_243 gnd vdd FILL
XFILL_13_BUFX4_13 gnd vdd FILL
XFILL_44_DFFSR_254 gnd vdd FILL
XFILL_3_NOR2X1_80 gnd vdd FILL
XFILL_13_BUFX4_24 gnd vdd FILL
XFILL_44_DFFSR_265 gnd vdd FILL
XFILL_2_CLKBUF1_30 gnd vdd FILL
XFILL_3_NOR2X1_91 gnd vdd FILL
XFILL_2_CLKBUF1_41 gnd vdd FILL
XFILL_13_BUFX4_35 gnd vdd FILL
XFILL_12_BUFX4_9 gnd vdd FILL
XFILL_10_MUX2X1_104 gnd vdd FILL
XFILL_13_BUFX4_46 gnd vdd FILL
XFILL_71_DFFSR_110 gnd vdd FILL
XFILL_54_4_1 gnd vdd FILL
XFILL_13_BUFX4_57 gnd vdd FILL
XFILL_10_MUX2X1_115 gnd vdd FILL
XFILL_71_DFFSR_121 gnd vdd FILL
XFILL_13_BUFX4_68 gnd vdd FILL
XFILL_10_MUX2X1_126 gnd vdd FILL
XFILL_48_DFFSR_220 gnd vdd FILL
XFILL_71_DFFSR_132 gnd vdd FILL
XFILL_48_DFFSR_231 gnd vdd FILL
XFILL_13_BUFX4_79 gnd vdd FILL
XFILL_71_DFFSR_143 gnd vdd FILL
XFILL_48_DFFSR_242 gnd vdd FILL
XFILL_10_MUX2X1_137 gnd vdd FILL
XFILL_71_DFFSR_154 gnd vdd FILL
XFILL_10_MUX2X1_148 gnd vdd FILL
XFILL_48_DFFSR_253 gnd vdd FILL
XFILL_71_DFFSR_165 gnd vdd FILL
XFILL_10_MUX2X1_159 gnd vdd FILL
XFILL_48_DFFSR_264 gnd vdd FILL
XFILL_71_DFFSR_176 gnd vdd FILL
XFILL_48_DFFSR_275 gnd vdd FILL
XFILL_7_NOR2X1_90 gnd vdd FILL
XFILL_71_DFFSR_187 gnd vdd FILL
XFILL_71_DFFSR_198 gnd vdd FILL
XFILL_75_DFFSR_120 gnd vdd FILL
XFILL_75_DFFSR_131 gnd vdd FILL
XFILL_11_OAI21X1_20 gnd vdd FILL
XFILL_11_OAI21X1_31 gnd vdd FILL
XFILL_0_DFFSR_1 gnd vdd FILL
XFILL_75_DFFSR_142 gnd vdd FILL
XFILL_11_OAI21X1_42 gnd vdd FILL
XFILL_75_DFFSR_153 gnd vdd FILL
XFILL_75_DFFSR_164 gnd vdd FILL
XFILL_75_DFFSR_175 gnd vdd FILL
XFILL_0_NOR2X1_170 gnd vdd FILL
XFILL_75_DFFSR_186 gnd vdd FILL
XFILL_0_NOR2X1_181 gnd vdd FILL
XFILL_75_DFFSR_197 gnd vdd FILL
XFILL_0_NOR2X1_192 gnd vdd FILL
XAOI22X1_9 INVX1_120/Y NOR2X1_19/A NOR2X1_16/A INVX1_121/Y gnd AOI22X1_9/Y vdd AOI22X1
XFILL_79_DFFSR_130 gnd vdd FILL
XFILL_79_DFFSR_141 gnd vdd FILL
XFILL_79_DFFSR_152 gnd vdd FILL
XFILL_7_INVX1_14 gnd vdd FILL
XFILL_79_DFFSR_163 gnd vdd FILL
XFILL_7_INVX1_25 gnd vdd FILL
XINVX1_208 DFFSR_77/Q gnd INVX1_208/Y vdd INVX1
XFILL_7_INVX1_36 gnd vdd FILL
XFILL_79_DFFSR_174 gnd vdd FILL
XFILL_79_DFFSR_185 gnd vdd FILL
XFILL_7_INVX1_47 gnd vdd FILL
XINVX1_219 DFFSR_71/Q gnd INVX1_219/Y vdd INVX1
XFILL_8_AND2X2_6 gnd vdd FILL
XFILL_79_DFFSR_196 gnd vdd FILL
XFILL_7_INVX1_58 gnd vdd FILL
XFILL_7_INVX1_69 gnd vdd FILL
XFILL_0_MUX2X1_110 gnd vdd FILL
XFILL_3_NAND2X1_2 gnd vdd FILL
XFILL_0_MUX2X1_121 gnd vdd FILL
XFILL_57_DFFSR_109 gnd vdd FILL
XFILL_0_MUX2X1_132 gnd vdd FILL
XFILL_35_DFFSR_3 gnd vdd FILL
XFILL_0_MUX2X1_143 gnd vdd FILL
XFILL_5_BUFX4_12 gnd vdd FILL
XFILL_5_BUFX4_23 gnd vdd FILL
XFILL_0_MUX2X1_154 gnd vdd FILL
XFILL_0_MUX2X1_165 gnd vdd FILL
XFILL_13_NAND3X1_18 gnd vdd FILL
XNAND2X1_19 BUFX4_58/Y NOR2X1_29/Y gnd OAI22X1_33/D vdd NAND2X1
XFILL_5_BUFX4_34 gnd vdd FILL
XFILL_5_BUFX4_45 gnd vdd FILL
XFILL_13_NAND3X1_29 gnd vdd FILL
XFILL_0_MUX2X1_176 gnd vdd FILL
XFILL_0_MUX2X1_187 gnd vdd FILL
XFILL_5_BUFX4_56 gnd vdd FILL
XFILL_7_NAND2X1_1 gnd vdd FILL
XFILL_5_BUFX4_67 gnd vdd FILL
XFILL_5_BUFX4_78 gnd vdd FILL
XFILL_33_CLKBUF1_18 gnd vdd FILL
XFILL_5_BUFX4_89 gnd vdd FILL
XFILL_11_DFFSR_210 gnd vdd FILL
XFILL_33_CLKBUF1_29 gnd vdd FILL
XFILL_11_DFFSR_221 gnd vdd FILL
XFILL_11_DFFSR_232 gnd vdd FILL
XFILL_11_DFFSR_243 gnd vdd FILL
XFILL_45_4_1 gnd vdd FILL
XFILL_11_DFFSR_254 gnd vdd FILL
XFILL_11_DFFSR_265 gnd vdd FILL
XFILL_15_DFFSR_220 gnd vdd FILL
XFILL_15_DFFSR_231 gnd vdd FILL
XFILL_15_DFFSR_242 gnd vdd FILL
XFILL_28_9 gnd vdd FILL
XFILL_15_DFFSR_253 gnd vdd FILL
XFILL_15_DFFSR_264 gnd vdd FILL
XFILL_15_DFFSR_275 gnd vdd FILL
XFILL_57_DFFSR_7 gnd vdd FILL
XFILL_42_DFFSR_120 gnd vdd FILL
XFILL_42_DFFSR_131 gnd vdd FILL
XFILL_3_AOI21X1_7 gnd vdd FILL
XFILL_19_DFFSR_230 gnd vdd FILL
XFILL_42_DFFSR_142 gnd vdd FILL
XFILL_19_DFFSR_241 gnd vdd FILL
XFILL_42_DFFSR_153 gnd vdd FILL
XFILL_19_DFFSR_252 gnd vdd FILL
XFILL_42_DFFSR_164 gnd vdd FILL
XFILL_42_DFFSR_175 gnd vdd FILL
XFILL_19_DFFSR_263 gnd vdd FILL
XFILL_19_DFFSR_274 gnd vdd FILL
XFILL_16_MUX2X1_19 gnd vdd FILL
XFILL_42_DFFSR_186 gnd vdd FILL
XFILL_42_DFFSR_197 gnd vdd FILL
XFILL_3_NAND3X1_13 gnd vdd FILL
XFILL_46_DFFSR_130 gnd vdd FILL
XFILL_7_AOI21X1_6 gnd vdd FILL
XFILL_3_NAND3X1_24 gnd vdd FILL
XFILL_3_NAND3X1_35 gnd vdd FILL
XFILL_46_DFFSR_141 gnd vdd FILL
XFILL_46_DFFSR_152 gnd vdd FILL
XFILL_3_NAND3X1_46 gnd vdd FILL
XNOR3X1_7 NOR3X1_7/A NOR3X1_7/B NOR3X1_7/C gnd NOR3X1_7/Y vdd NOR3X1
XFILL_3_NAND3X1_57 gnd vdd FILL
XFILL_46_DFFSR_163 gnd vdd FILL
XFILL_46_DFFSR_174 gnd vdd FILL
XFILL_3_NAND3X1_68 gnd vdd FILL
XFILL_7_NAND2X1_15 gnd vdd FILL
XFILL_7_NAND2X1_26 gnd vdd FILL
XFILL_46_DFFSR_185 gnd vdd FILL
XFILL_3_NAND3X1_79 gnd vdd FILL
XFILL_7_NAND2X1_37 gnd vdd FILL
XFILL_7_NAND2X1_48 gnd vdd FILL
XFILL_46_DFFSR_196 gnd vdd FILL
XFILL_7_NAND2X1_59 gnd vdd FILL
XFILL_12_AOI22X1_3 gnd vdd FILL
XFILL_5_1 gnd vdd FILL
XFILL_24_DFFSR_109 gnd vdd FILL
XFILL_17_MUX2X1_190 gnd vdd FILL
XFILL_61_3 gnd vdd FILL
XFILL_16_AOI22X1_2 gnd vdd FILL
XFILL_54_2 gnd vdd FILL
XFILL_1_DFFSR_19 gnd vdd FILL
XFILL_28_DFFSR_108 gnd vdd FILL
XFILL_11_NOR2X1_7 gnd vdd FILL
XFILL_28_DFFSR_119 gnd vdd FILL
XFILL_36_4_1 gnd vdd FILL
XFILL_3_INVX1_40 gnd vdd FILL
XFILL_3_INVX1_51 gnd vdd FILL
XFILL_3_INVX1_62 gnd vdd FILL
XFILL_3_INVX1_73 gnd vdd FILL
XFILL_49_DFFSR_10 gnd vdd FILL
XFILL_49_DFFSR_21 gnd vdd FILL
XFILL_3_INVX1_84 gnd vdd FILL
XFILL_3_INVX1_95 gnd vdd FILL
XFILL_49_DFFSR_32 gnd vdd FILL
XFILL_49_DFFSR_43 gnd vdd FILL
XFILL_49_DFFSR_54 gnd vdd FILL
XFILL_49_DFFSR_65 gnd vdd FILL
XFILL_10_MUX2X1_5 gnd vdd FILL
XFILL_49_DFFSR_76 gnd vdd FILL
XFILL_49_DFFSR_87 gnd vdd FILL
XFILL_49_DFFSR_98 gnd vdd FILL
XFILL_22_CLKBUF1_14 gnd vdd FILL
XFILL_22_CLKBUF1_25 gnd vdd FILL
XFILL_22_CLKBUF1_36 gnd vdd FILL
XFILL_74_DFFSR_209 gnd vdd FILL
XFILL_1_BUFX4_60 gnd vdd FILL
XFILL_18_DFFSR_20 gnd vdd FILL
XFILL_18_DFFSR_31 gnd vdd FILL
XFILL_1_BUFX4_71 gnd vdd FILL
XFILL_18_DFFSR_42 gnd vdd FILL
XFILL_5_CLKBUF1_18 gnd vdd FILL
XFILL_18_DFFSR_53 gnd vdd FILL
XFILL_1_BUFX4_82 gnd vdd FILL
XFILL_28_NOR3X1_19 gnd vdd FILL
XFILL_5_CLKBUF1_29 gnd vdd FILL
XFILL_1_BUFX4_93 gnd vdd FILL
XFILL_18_DFFSR_64 gnd vdd FILL
XFILL_18_DFFSR_75 gnd vdd FILL
XFILL_13_DFFSR_130 gnd vdd FILL
XFILL_78_DFFSR_208 gnd vdd FILL
XFILL_18_DFFSR_86 gnd vdd FILL
XFILL_0_AOI21X1_15 gnd vdd FILL
XFILL_78_DFFSR_219 gnd vdd FILL
XFILL_0_AOI21X1_26 gnd vdd FILL
XFILL_18_DFFSR_97 gnd vdd FILL
XFILL_0_AOI21X1_37 gnd vdd FILL
XFILL_13_DFFSR_141 gnd vdd FILL
XFILL_13_DFFSR_152 gnd vdd FILL
XFILL_0_AOI21X1_48 gnd vdd FILL
XFILL_58_DFFSR_30 gnd vdd FILL
XFILL_13_DFFSR_163 gnd vdd FILL
XFILL_0_AOI21X1_59 gnd vdd FILL
XFILL_13_DFFSR_174 gnd vdd FILL
XFILL_10_OAI22X1_17 gnd vdd FILL
XFILL_58_DFFSR_41 gnd vdd FILL
XFILL_29_NOR3X1_5 gnd vdd FILL
XFILL_10_OAI22X1_28 gnd vdd FILL
XFILL_58_DFFSR_52 gnd vdd FILL
XFILL_2_CLKBUF1_6 gnd vdd FILL
XFILL_58_DFFSR_63 gnd vdd FILL
XFILL_13_DFFSR_185 gnd vdd FILL
XFILL_10_OAI22X1_39 gnd vdd FILL
XFILL_13_DFFSR_196 gnd vdd FILL
XFILL_3_NOR2X1_103 gnd vdd FILL
XFILL_58_DFFSR_74 gnd vdd FILL
XFILL_58_DFFSR_85 gnd vdd FILL
XFILL_3_NOR2X1_114 gnd vdd FILL
XFILL_3_NOR2X1_125 gnd vdd FILL
XFILL_17_DFFSR_140 gnd vdd FILL
XFILL_14_OAI21X1_19 gnd vdd FILL
XFILL_58_DFFSR_96 gnd vdd FILL
XFILL_4_DFFSR_2 gnd vdd FILL
XFILL_3_NOR2X1_136 gnd vdd FILL
XFILL_17_DFFSR_151 gnd vdd FILL
XFILL_17_DFFSR_162 gnd vdd FILL
XFILL_3_NOR2X1_147 gnd vdd FILL
XFILL_3_NOR2X1_6 gnd vdd FILL
XFILL_3_NOR2X1_158 gnd vdd FILL
XFILL_17_DFFSR_173 gnd vdd FILL
XFILL_74_DFFSR_1 gnd vdd FILL
XFILL_6_CLKBUF1_5 gnd vdd FILL
XFILL_17_DFFSR_184 gnd vdd FILL
XFILL_3_NOR2X1_169 gnd vdd FILL
XFILL_17_DFFSR_195 gnd vdd FILL
XFILL_27_DFFSR_40 gnd vdd FILL
XFILL_27_DFFSR_51 gnd vdd FILL
XFILL_27_DFFSR_62 gnd vdd FILL
XFILL_27_DFFSR_73 gnd vdd FILL
XFILL_2_BUFX4_100 gnd vdd FILL
XFILL_27_DFFSR_84 gnd vdd FILL
XFILL_27_DFFSR_95 gnd vdd FILL
XFILL_27_4_1 gnd vdd FILL
XFILL_2_4_1 gnd vdd FILL
XFILL_13_NOR3X1_30 gnd vdd FILL
XFILL_13_NOR3X1_41 gnd vdd FILL
XFILL_13_NOR3X1_52 gnd vdd FILL
XFILL_2_MUX2X1_4 gnd vdd FILL
XFILL_20_MUX2X1_105 gnd vdd FILL
XFILL_20_MUX2X1_116 gnd vdd FILL
XFILL_67_DFFSR_50 gnd vdd FILL
XFILL_20_MUX2X1_127 gnd vdd FILL
XFILL_67_DFFSR_61 gnd vdd FILL
XFILL_63_DFFSR_230 gnd vdd FILL
XFILL_67_DFFSR_72 gnd vdd FILL
XFILL_67_DFFSR_83 gnd vdd FILL
XFILL_63_DFFSR_241 gnd vdd FILL
XFILL_20_MUX2X1_138 gnd vdd FILL
XFILL_20_MUX2X1_149 gnd vdd FILL
XFILL_63_DFFSR_252 gnd vdd FILL
XFILL_67_DFFSR_94 gnd vdd FILL
XFILL_63_DFFSR_263 gnd vdd FILL
XFILL_63_DFFSR_274 gnd vdd FILL
XFILL_3_MUX2X1_109 gnd vdd FILL
XFILL_17_NOR3X1_40 gnd vdd FILL
XFILL_39_DFFSR_4 gnd vdd FILL
XFILL_17_NOR3X1_51 gnd vdd FILL
XFILL_8_NOR2X1_203 gnd vdd FILL
XFILL_0_OAI22X1_12 gnd vdd FILL
XFILL_0_OAI22X1_23 gnd vdd FILL
XFILL_67_DFFSR_240 gnd vdd FILL
XFILL_67_DFFSR_251 gnd vdd FILL
XFILL_0_OAI22X1_34 gnd vdd FILL
XFILL_67_DFFSR_262 gnd vdd FILL
XFILL_10_3_1 gnd vdd FILL
XFILL_0_OAI22X1_45 gnd vdd FILL
XFILL_22_CLKBUF1_3 gnd vdd FILL
XFILL_36_DFFSR_60 gnd vdd FILL
XFILL_4_OAI21X1_14 gnd vdd FILL
XFILL_67_DFFSR_273 gnd vdd FILL
XFILL_36_DFFSR_71 gnd vdd FILL
XFILL_36_DFFSR_82 gnd vdd FILL
XFILL_4_OAI21X1_25 gnd vdd FILL
XFILL_36_DFFSR_93 gnd vdd FILL
XFILL_0_NOR2X1_13 gnd vdd FILL
XFILL_4_OAI21X1_36 gnd vdd FILL
XFILL_0_NOR2X1_24 gnd vdd FILL
XFILL_41_DFFSR_209 gnd vdd FILL
XFILL_0_NOR2X1_35 gnd vdd FILL
XFILL_4_OAI21X1_47 gnd vdd FILL
XAOI21X1_50 MUX2X1_8/A NOR2X1_9/B NOR2X1_8/Y gnd DFFSR_267/D vdd AOI21X1
XFILL_0_NOR2X1_46 gnd vdd FILL
XAOI21X1_61 OAI21X1_42/Y NAND3X1_43/B NAND3X1_43/A gnd AND2X2_1/B vdd AOI21X1
XFILL_0_NOR2X1_57 gnd vdd FILL
XAOI21X1_72 DFFSR_151/Q NOR2X1_43/Y NOR2X1_98/Y gnd NAND3X1_10/B vdd AOI21X1
XFILL_0_NOR2X1_68 gnd vdd FILL
XFILL_0_NOR2X1_79 gnd vdd FILL
XFILL_26_CLKBUF1_2 gnd vdd FILL
XFILL_76_DFFSR_70 gnd vdd FILL
XFILL_76_DFFSR_81 gnd vdd FILL
XFILL_76_DFFSR_92 gnd vdd FILL
XOAI21X1_1 OAI21X1_1/A OAI21X1_1/B OAI21X1_1/C gnd OAI21X1_1/Y vdd OAI21X1
XFILL_4_NOR2X1_12 gnd vdd FILL
XFILL_45_DFFSR_208 gnd vdd FILL
XFILL_4_NOR2X1_23 gnd vdd FILL
XFILL_45_DFFSR_219 gnd vdd FILL
XFILL_4_NOR2X1_34 gnd vdd FILL
XFILL_7_OAI21X1_9 gnd vdd FILL
XFILL_3_NAND2X1_90 gnd vdd FILL
XFILL_4_NOR2X1_45 gnd vdd FILL
XFILL_4_NOR2X1_56 gnd vdd FILL
XFILL_9_0_0 gnd vdd FILL
XFILL_4_NOR2X1_67 gnd vdd FILL
XFILL_4_NOR2X1_78 gnd vdd FILL
XFILL_4_NOR2X1_89 gnd vdd FILL
XFILL_11_CLKBUF1_10 gnd vdd FILL
XFILL_49_DFFSR_207 gnd vdd FILL
XFILL_11_CLKBUF1_21 gnd vdd FILL
XFILL_72_DFFSR_108 gnd vdd FILL
XFILL_8_NOR2X1_11 gnd vdd FILL
XFILL_11_CLKBUF1_32 gnd vdd FILL
XFILL_72_DFFSR_119 gnd vdd FILL
XFILL_8_NOR2X1_22 gnd vdd FILL
XFILL_8_NOR2X1_33 gnd vdd FILL
XFILL_49_DFFSR_218 gnd vdd FILL
XFILL_8_NOR2X1_44 gnd vdd FILL
XFILL_49_DFFSR_229 gnd vdd FILL
XFILL_45_DFFSR_80 gnd vdd FILL
XFILL_8_NOR2X1_55 gnd vdd FILL
XFILL_12_OAI22X1_6 gnd vdd FILL
XFILL_45_DFFSR_91 gnd vdd FILL
XFILL_8_NOR2X1_66 gnd vdd FILL
XFILL_8_NOR2X1_77 gnd vdd FILL
XFILL_8_NOR2X1_88 gnd vdd FILL
XFILL_8_NOR2X1_99 gnd vdd FILL
XFILL_76_DFFSR_107 gnd vdd FILL
XFILL_76_DFFSR_118 gnd vdd FILL
XFILL_76_DFFSR_129 gnd vdd FILL
XFILL_18_4_1 gnd vdd FILL
XFILL_85_DFFSR_90 gnd vdd FILL
XFILL_16_OAI22X1_5 gnd vdd FILL
XFILL_61_7_2 gnd vdd FILL
XFILL_14_DFFSR_90 gnd vdd FILL
XFILL_60_2_1 gnd vdd FILL
XFILL_26_6 gnd vdd FILL
XFILL_30_DFFSR_230 gnd vdd FILL
XFILL_30_DFFSR_241 gnd vdd FILL
XFILL_30_DFFSR_252 gnd vdd FILL
XFILL_19_5 gnd vdd FILL
XFILL_30_DFFSR_263 gnd vdd FILL
XFILL_30_DFFSR_274 gnd vdd FILL
XFILL_34_DFFSR_240 gnd vdd FILL
XFILL_34_DFFSR_251 gnd vdd FILL
XFILL_34_DFFSR_262 gnd vdd FILL
XFILL_34_DFFSR_273 gnd vdd FILL
XFILL_0_MUX2X1_20 gnd vdd FILL
XFILL_0_MUX2X1_31 gnd vdd FILL
XFILL_0_MUX2X1_42 gnd vdd FILL
XFILL_0_MUX2X1_53 gnd vdd FILL
XFILL_0_MUX2X1_64 gnd vdd FILL
XFILL_61_DFFSR_140 gnd vdd FILL
XFILL_0_MUX2X1_75 gnd vdd FILL
XFILL_0_MUX2X1_86 gnd vdd FILL
XFILL_61_DFFSR_151 gnd vdd FILL
XFILL_38_DFFSR_250 gnd vdd FILL
XFILL_61_DFFSR_162 gnd vdd FILL
XFILL_38_DFFSR_261 gnd vdd FILL
XFILL_0_MUX2X1_97 gnd vdd FILL
XFILL_61_DFFSR_173 gnd vdd FILL
XFILL_61_DFFSR_184 gnd vdd FILL
XFILL_38_DFFSR_272 gnd vdd FILL
XFILL_4_MUX2X1_30 gnd vdd FILL
XFILL_61_DFFSR_195 gnd vdd FILL
XFILL_4_MUX2X1_41 gnd vdd FILL
XFILL_12_DFFSR_208 gnd vdd FILL
XFILL_12_DFFSR_219 gnd vdd FILL
XFILL_4_MUX2X1_52 gnd vdd FILL
XFILL_4_MUX2X1_63 gnd vdd FILL
XFILL_4_MUX2X1_74 gnd vdd FILL
XFILL_4_MUX2X1_85 gnd vdd FILL
XFILL_10_OAI21X1_50 gnd vdd FILL
XFILL_65_DFFSR_150 gnd vdd FILL
XFILL_65_DFFSR_161 gnd vdd FILL
XFILL_4_MUX2X1_96 gnd vdd FILL
XFILL_65_DFFSR_172 gnd vdd FILL
XFILL_65_DFFSR_183 gnd vdd FILL
XFILL_65_DFFSR_194 gnd vdd FILL
XFILL_10_BUFX4_17 gnd vdd FILL
XFILL_8_MUX2X1_40 gnd vdd FILL
XFILL_16_DFFSR_207 gnd vdd FILL
XFILL_10_BUFX4_28 gnd vdd FILL
XFILL_8_MUX2X1_51 gnd vdd FILL
XFILL_13_NAND3X1_7 gnd vdd FILL
XFILL_16_DFFSR_218 gnd vdd FILL
XFILL_8_MUX2X1_62 gnd vdd FILL
XFILL_10_BUFX4_39 gnd vdd FILL
XFILL_16_DFFSR_229 gnd vdd FILL
XFILL_8_MUX2X1_73 gnd vdd FILL
XFILL_8_MUX2X1_84 gnd vdd FILL
XFILL_69_DFFSR_160 gnd vdd FILL
XFILL_8_MUX2X1_95 gnd vdd FILL
XFILL_69_DFFSR_171 gnd vdd FILL
XFILL_69_DFFSR_182 gnd vdd FILL
XFILL_69_DFFSR_193 gnd vdd FILL
XFILL_43_DFFSR_107 gnd vdd FILL
XFILL_43_DFFSR_118 gnd vdd FILL
XFILL_43_DFFSR_129 gnd vdd FILL
XFILL_52_7_2 gnd vdd FILL
XFILL_51_2_1 gnd vdd FILL
XFILL_47_DFFSR_106 gnd vdd FILL
XFILL_40_DFFSR_4 gnd vdd FILL
XFILL_47_DFFSR_117 gnd vdd FILL
XFILL_8_DFFSR_3 gnd vdd FILL
XFILL_47_DFFSR_128 gnd vdd FILL
XFILL_47_DFFSR_139 gnd vdd FILL
XFILL_20_MUX2X1_50 gnd vdd FILL
XFILL_12_NAND3X1_15 gnd vdd FILL
XFILL_20_MUX2X1_61 gnd vdd FILL
XFILL_12_NAND3X1_26 gnd vdd FILL
XFILL_20_MUX2X1_72 gnd vdd FILL
XFILL_20_MUX2X1_83 gnd vdd FILL
XFILL_12_NAND3X1_37 gnd vdd FILL
XFILL_78_DFFSR_2 gnd vdd FILL
XFILL_12_NAND3X1_48 gnd vdd FILL
XFILL_12_NAND3X1_59 gnd vdd FILL
XFILL_20_MUX2X1_94 gnd vdd FILL
XFILL_4_INVX1_18 gnd vdd FILL
XFILL_4_INVX1_29 gnd vdd FILL
XFILL_32_CLKBUF1_15 gnd vdd FILL
XFILL_32_CLKBUF1_26 gnd vdd FILL
XFILL_32_CLKBUF1_37 gnd vdd FILL
XFILL_3_BUFX2_9 gnd vdd FILL
XFILL_2_BUFX4_16 gnd vdd FILL
XFILL_2_BUFX4_27 gnd vdd FILL
XFILL_62_DFFSR_8 gnd vdd FILL
XFILL_2_BUFX4_38 gnd vdd FILL
XFILL_2_BUFX4_49 gnd vdd FILL
XFILL_59_3_1 gnd vdd FILL
XFILL_32_DFFSR_150 gnd vdd FILL
XFILL_32_DFFSR_161 gnd vdd FILL
XFILL_32_DFFSR_172 gnd vdd FILL
XFILL_32_DFFSR_183 gnd vdd FILL
XFILL_59_DFFSR_19 gnd vdd FILL
XFILL_32_DFFSR_194 gnd vdd FILL
XFILL_2_NAND3X1_10 gnd vdd FILL
XFILL_2_NAND3X1_21 gnd vdd FILL
XFILL_2_NAND3X1_32 gnd vdd FILL
XFILL_2_NAND3X1_43 gnd vdd FILL
XFILL_36_DFFSR_160 gnd vdd FILL
XFILL_2_NAND3X1_54 gnd vdd FILL
XFILL_2_NAND3X1_65 gnd vdd FILL
XFILL_6_NAND2X1_12 gnd vdd FILL
XFILL_36_DFFSR_171 gnd vdd FILL
XFILL_6_NAND2X1_23 gnd vdd FILL
XFILL_2_NAND3X1_76 gnd vdd FILL
XFILL_36_DFFSR_182 gnd vdd FILL
XFILL_36_DFFSR_193 gnd vdd FILL
XFILL_6_NAND2X1_34 gnd vdd FILL
XFILL_10_DFFSR_107 gnd vdd FILL
XFILL_2_BUFX4_3 gnd vdd FILL
XFILL_43_7_2 gnd vdd FILL
XFILL_2_NAND3X1_87 gnd vdd FILL
XFILL_6_NAND2X1_45 gnd vdd FILL
XFILL_10_DFFSR_118 gnd vdd FILL
XFILL_6_NAND2X1_56 gnd vdd FILL
XFILL_2_NAND3X1_98 gnd vdd FILL
XFILL_15_BUFX4_1 gnd vdd FILL
XFILL_42_2_1 gnd vdd FILL
XFILL_10_DFFSR_129 gnd vdd FILL
XFILL_6_NAND2X1_67 gnd vdd FILL
XFILL_6_NAND2X1_78 gnd vdd FILL
XMUX2X1_5 MUX2X1_5/A MUX2X1_9/A MUX2X1_7/S gnd MUX2X1_5/Y vdd MUX2X1
XFILL_28_DFFSR_18 gnd vdd FILL
XFILL_6_NAND2X1_89 gnd vdd FILL
XFILL_28_DFFSR_29 gnd vdd FILL
XFILL_14_DFFSR_106 gnd vdd FILL
XFILL_14_DFFSR_117 gnd vdd FILL
XFILL_14_DFFSR_128 gnd vdd FILL
XFILL_68_DFFSR_17 gnd vdd FILL
XFILL_14_DFFSR_139 gnd vdd FILL
XFILL_68_DFFSR_28 gnd vdd FILL
XFILL_68_DFFSR_39 gnd vdd FILL
XFILL_82_DFFSR_250 gnd vdd FILL
XFILL_82_DFFSR_261 gnd vdd FILL
XFILL_18_DFFSR_105 gnd vdd FILL
XFILL_82_DFFSR_272 gnd vdd FILL
XFILL_18_DFFSR_116 gnd vdd FILL
XFILL_18_DFFSR_127 gnd vdd FILL
XFILL_1_INVX1_7 gnd vdd FILL
XFILL_18_DFFSR_138 gnd vdd FILL
XFILL_18_DFFSR_149 gnd vdd FILL
XFILL_13_AOI21X1_1 gnd vdd FILL
XCLKBUF1_6 BUFX4_95/Y gnd CLKBUF1_6/Y vdd CLKBUF1
XFILL_6_AOI22X1_10 gnd vdd FILL
XFILL_86_DFFSR_260 gnd vdd FILL
XFILL_10_NOR3X1_18 gnd vdd FILL
XFILL_37_DFFSR_16 gnd vdd FILL
XFILL_86_DFFSR_271 gnd vdd FILL
XFILL_37_DFFSR_27 gnd vdd FILL
XFILL_10_NOR3X1_29 gnd vdd FILL
XFILL_37_DFFSR_38 gnd vdd FILL
XFILL_60_DFFSR_207 gnd vdd FILL
XFILL_37_DFFSR_49 gnd vdd FILL
XFILL_60_DFFSR_218 gnd vdd FILL
XFILL_60_DFFSR_229 gnd vdd FILL
XFILL_14_NOR3X1_17 gnd vdd FILL
XFILL_77_DFFSR_15 gnd vdd FILL
XFILL_14_NOR3X1_28 gnd vdd FILL
XFILL_77_DFFSR_26 gnd vdd FILL
XFILL_21_CLKBUF1_11 gnd vdd FILL
XFILL_77_DFFSR_37 gnd vdd FILL
XFILL_14_NOR3X1_39 gnd vdd FILL
XFILL_21_CLKBUF1_22 gnd vdd FILL
XFILL_64_DFFSR_206 gnd vdd FILL
XFILL_21_CLKBUF1_33 gnd vdd FILL
XFILL_77_DFFSR_48 gnd vdd FILL
XBUFX4_100 INVX8_3/Y gnd MUX2X1_2/A vdd BUFX4
XFILL_64_DFFSR_217 gnd vdd FILL
XFILL_77_DFFSR_59 gnd vdd FILL
XFILL_64_DFFSR_228 gnd vdd FILL
XFILL_64_DFFSR_239 gnd vdd FILL
XFILL_0_INVX1_11 gnd vdd FILL
XFILL_0_INVX1_22 gnd vdd FILL
XFILL_18_NOR3X1_16 gnd vdd FILL
XFILL_4_CLKBUF1_15 gnd vdd FILL
XFILL_0_INVX1_33 gnd vdd FILL
XFILL_18_NOR3X1_27 gnd vdd FILL
XFILL_4_CLKBUF1_26 gnd vdd FILL
XFILL_0_INVX1_44 gnd vdd FILL
XFILL_1_AND2X2_3 gnd vdd FILL
XFILL_5_INVX8_1 gnd vdd FILL
XFILL_18_NOR3X1_38 gnd vdd FILL
XFILL_0_INVX1_55 gnd vdd FILL
XFILL_4_CLKBUF1_37 gnd vdd FILL
XNOR2X1_204 DFFSR_275/Q MUX2X1_22/S gnd NOR2X1_204/Y vdd NOR2X1
XFILL_18_NOR3X1_49 gnd vdd FILL
XFILL_68_DFFSR_205 gnd vdd FILL
XFILL_0_INVX1_66 gnd vdd FILL
XFILL_0_INVX1_77 gnd vdd FILL
XFILL_68_DFFSR_216 gnd vdd FILL
XFILL_46_DFFSR_14 gnd vdd FILL
XFILL_0_INVX1_88 gnd vdd FILL
XFILL_68_DFFSR_227 gnd vdd FILL
XFILL_46_DFFSR_25 gnd vdd FILL
XFILL_0_INVX1_99 gnd vdd FILL
XFILL_46_DFFSR_36 gnd vdd FILL
XFILL_34_7_2 gnd vdd FILL
XFILL_68_DFFSR_238 gnd vdd FILL
XFILL_68_DFFSR_249 gnd vdd FILL
XFILL_31_4 gnd vdd FILL
XFILL_46_DFFSR_47 gnd vdd FILL
XFILL_46_DFFSR_58 gnd vdd FILL
XFILL_33_2_1 gnd vdd FILL
XFILL_46_DFFSR_69 gnd vdd FILL
XFILL_24_3 gnd vdd FILL
XFILL_2_NOR2X1_100 gnd vdd FILL
XFILL_13_OAI21X1_16 gnd vdd FILL
XFILL_2_NOR2X1_111 gnd vdd FILL
XFILL_86_DFFSR_13 gnd vdd FILL
XFILL_2_NOR2X1_122 gnd vdd FILL
XFILL_13_OAI21X1_27 gnd vdd FILL
XFILL_86_DFFSR_24 gnd vdd FILL
XFILL_2_NOR2X1_133 gnd vdd FILL
XFILL_86_DFFSR_35 gnd vdd FILL
XFILL_2_NOR2X1_144 gnd vdd FILL
XFILL_13_OAI21X1_38 gnd vdd FILL
XFILL_22_DFFSR_1 gnd vdd FILL
XFILL_17_2 gnd vdd FILL
XFILL_13_OAI21X1_49 gnd vdd FILL
XFILL_86_DFFSR_46 gnd vdd FILL
XFILL_86_DFFSR_57 gnd vdd FILL
XFILL_2_NOR2X1_155 gnd vdd FILL
XFILL_15_DFFSR_13 gnd vdd FILL
XFILL_2_NOR2X1_166 gnd vdd FILL
XFILL_86_DFFSR_68 gnd vdd FILL
XFILL_15_DFFSR_24 gnd vdd FILL
XFILL_2_NOR2X1_177 gnd vdd FILL
XFILL_15_DFFSR_35 gnd vdd FILL
XFILL_2_NOR2X1_188 gnd vdd FILL
XFILL_86_DFFSR_79 gnd vdd FILL
XFILL_15_DFFSR_46 gnd vdd FILL
XFILL_15_DFFSR_57 gnd vdd FILL
XFILL_2_NOR2X1_199 gnd vdd FILL
XFILL_26_13 gnd vdd FILL
XFILL_15_DFFSR_68 gnd vdd FILL
XFILL_15_DFFSR_79 gnd vdd FILL
XFILL_55_DFFSR_12 gnd vdd FILL
XFILL_55_DFFSR_23 gnd vdd FILL
XFILL_55_DFFSR_34 gnd vdd FILL
XFILL_26_NOR3X1_9 gnd vdd FILL
XFILL_55_DFFSR_45 gnd vdd FILL
XFILL_55_DFFSR_56 gnd vdd FILL
XFILL_55_DFFSR_67 gnd vdd FILL
XFILL_55_DFFSR_78 gnd vdd FILL
XFILL_55_DFFSR_89 gnd vdd FILL
XFILL_53_DFFSR_260 gnd vdd FILL
XFILL_2_MUX2X1_106 gnd vdd FILL
XFILL_53_DFFSR_271 gnd vdd FILL
XFILL_2_MUX2X1_117 gnd vdd FILL
XFILL_44_DFFSR_5 gnd vdd FILL
XFILL_24_DFFSR_11 gnd vdd FILL
XFILL_2_MUX2X1_128 gnd vdd FILL
XFILL_7_NOR2X1_200 gnd vdd FILL
XFILL_24_DFFSR_22 gnd vdd FILL
XFILL_2_MUX2X1_139 gnd vdd FILL
XFILL_24_DFFSR_33 gnd vdd FILL
XFILL_24_DFFSR_44 gnd vdd FILL
XFILL_24_DFFSR_55 gnd vdd FILL
XFILL_80_DFFSR_160 gnd vdd FILL
XFILL_24_DFFSR_66 gnd vdd FILL
XFILL_24_DFFSR_77 gnd vdd FILL
XFILL_80_DFFSR_171 gnd vdd FILL
XFILL_3_OAI21X1_11 gnd vdd FILL
XFILL_57_DFFSR_270 gnd vdd FILL
XFILL_80_DFFSR_182 gnd vdd FILL
XFILL_24_DFFSR_88 gnd vdd FILL
XFILL_3_OAI21X1_22 gnd vdd FILL
XFILL_24_DFFSR_99 gnd vdd FILL
XFILL_80_DFFSR_193 gnd vdd FILL
XFILL_3_OAI21X1_33 gnd vdd FILL
XFILL_64_DFFSR_10 gnd vdd FILL
XFILL_31_DFFSR_206 gnd vdd FILL
XFILL_64_DFFSR_21 gnd vdd FILL
XFILL_31_DFFSR_217 gnd vdd FILL
XFILL_0_DFFSR_230 gnd vdd FILL
XFILL_64_DFFSR_32 gnd vdd FILL
XFILL_3_OAI21X1_44 gnd vdd FILL
XFILL_0_DFFSR_241 gnd vdd FILL
XFILL_31_DFFSR_228 gnd vdd FILL
XFILL_64_DFFSR_43 gnd vdd FILL
XFILL_31_DFFSR_239 gnd vdd FILL
XFILL_0_DFFSR_252 gnd vdd FILL
XFILL_64_DFFSR_54 gnd vdd FILL
XFILL_64_DFFSR_65 gnd vdd FILL
XFILL_0_DFFSR_263 gnd vdd FILL
XFILL_64_DFFSR_76 gnd vdd FILL
XFILL_0_DFFSR_274 gnd vdd FILL
XFILL_84_DFFSR_170 gnd vdd FILL
XFILL_64_DFFSR_87 gnd vdd FILL
XFILL_84_DFFSR_181 gnd vdd FILL
XFILL_84_DFFSR_192 gnd vdd FILL
XFILL_35_DFFSR_205 gnd vdd FILL
XFILL_64_DFFSR_98 gnd vdd FILL
XFILL_25_7_2 gnd vdd FILL
XFILL_0_7_2 gnd vdd FILL
XFILL_7_DFFSR_12 gnd vdd FILL
XFILL_35_DFFSR_216 gnd vdd FILL
XFILL_35_DFFSR_227 gnd vdd FILL
XFILL_4_DFFSR_240 gnd vdd FILL
XFILL_7_DFFSR_23 gnd vdd FILL
XFILL_24_2_1 gnd vdd FILL
XFILL_4_DFFSR_251 gnd vdd FILL
XFILL_35_DFFSR_238 gnd vdd FILL
XFILL_35_DFFSR_249 gnd vdd FILL
XFILL_4_DFFSR_262 gnd vdd FILL
XFILL_7_DFFSR_34 gnd vdd FILL
XFILL_66_DFFSR_9 gnd vdd FILL
XFILL_33_DFFSR_20 gnd vdd FILL
XFILL_7_DFFSR_45 gnd vdd FILL
XFILL_7_DFFSR_56 gnd vdd FILL
XFILL_4_DFFSR_273 gnd vdd FILL
XFILL_33_DFFSR_31 gnd vdd FILL
XFILL_7_DFFSR_67 gnd vdd FILL
XFILL_1_MUX2X1_18 gnd vdd FILL
XFILL_33_DFFSR_42 gnd vdd FILL
XFILL_7_DFFSR_78 gnd vdd FILL
XFILL_1_MUX2X1_29 gnd vdd FILL
XFILL_62_DFFSR_105 gnd vdd FILL
XFILL_33_DFFSR_53 gnd vdd FILL
XFILL_39_DFFSR_204 gnd vdd FILL
XFILL_7_DFFSR_89 gnd vdd FILL
XFILL_39_DFFSR_215 gnd vdd FILL
XFILL_62_DFFSR_116 gnd vdd FILL
XFILL_33_DFFSR_64 gnd vdd FILL
XFILL_62_DFFSR_127 gnd vdd FILL
XFILL_10_CLKBUF1_40 gnd vdd FILL
XFILL_33_DFFSR_75 gnd vdd FILL
XFILL_33_DFFSR_86 gnd vdd FILL
XFILL_39_DFFSR_226 gnd vdd FILL
XFILL_62_DFFSR_138 gnd vdd FILL
XFILL_39_DFFSR_237 gnd vdd FILL
XFILL_8_DFFSR_250 gnd vdd FILL
XFILL_33_DFFSR_97 gnd vdd FILL
XFILL_62_DFFSR_149 gnd vdd FILL
XFILL_39_DFFSR_248 gnd vdd FILL
XFILL_8_DFFSR_261 gnd vdd FILL
XFILL_39_DFFSR_259 gnd vdd FILL
XFILL_8_DFFSR_272 gnd vdd FILL
XFILL_73_DFFSR_30 gnd vdd FILL
XFILL_73_DFFSR_41 gnd vdd FILL
XFILL_5_MUX2X1_17 gnd vdd FILL
XFILL_73_DFFSR_52 gnd vdd FILL
XFILL_5_MUX2X1_28 gnd vdd FILL
XFILL_66_DFFSR_104 gnd vdd FILL
XFILL_5_MUX2X1_39 gnd vdd FILL
XFILL_73_DFFSR_63 gnd vdd FILL
XFILL_66_DFFSR_115 gnd vdd FILL
XFILL_73_DFFSR_74 gnd vdd FILL
XFILL_66_DFFSR_126 gnd vdd FILL
XFILL_66_DFFSR_137 gnd vdd FILL
XFILL_73_DFFSR_85 gnd vdd FILL
XFILL_73_DFFSR_96 gnd vdd FILL
XFILL_66_DFFSR_148 gnd vdd FILL
XFILL_66_DFFSR_159 gnd vdd FILL
XFILL_9_MUX2X1_16 gnd vdd FILL
XFILL_6_BUFX4_4 gnd vdd FILL
XFILL_9_MUX2X1_27 gnd vdd FILL
XFILL_9_MUX2X1_38 gnd vdd FILL
XFILL_9_MUX2X1_49 gnd vdd FILL
XFILL_42_DFFSR_40 gnd vdd FILL
XFILL_1_AOI22X1_1 gnd vdd FILL
XFILL_13_NOR3X1_4 gnd vdd FILL
XFILL_19_MUX2X1_120 gnd vdd FILL
XFILL_42_DFFSR_51 gnd vdd FILL
XFILL_13_OAI21X1_4 gnd vdd FILL
XFILL_42_DFFSR_62 gnd vdd FILL
XFILL_19_MUX2X1_131 gnd vdd FILL
XFILL_10_NOR2X1_40 gnd vdd FILL
XFILL_19_MUX2X1_142 gnd vdd FILL
XFILL_10_NOR2X1_51 gnd vdd FILL
XFILL_42_DFFSR_73 gnd vdd FILL
XFILL_42_DFFSR_84 gnd vdd FILL
XFILL_19_MUX2X1_153 gnd vdd FILL
XFILL_10_NOR2X1_62 gnd vdd FILL
XFILL_20_DFFSR_260 gnd vdd FILL
XFILL_42_DFFSR_95 gnd vdd FILL
XFILL_20_DFFSR_271 gnd vdd FILL
XFILL_1_INVX1_200 gnd vdd FILL
XFILL_19_MUX2X1_164 gnd vdd FILL
XFILL_7_3_1 gnd vdd FILL
XFILL_10_NOR2X1_73 gnd vdd FILL
XFILL_19_MUX2X1_175 gnd vdd FILL
XBUFX4_17 BUFX4_47/A gnd DFFSR_89/R vdd BUFX4
XFILL_10_NOR2X1_84 gnd vdd FILL
XBUFX4_28 BUFX4_3/Y gnd DFFSR_64/R vdd BUFX4
XFILL_10_NOR2X1_95 gnd vdd FILL
XFILL_19_MUX2X1_186 gnd vdd FILL
XFILL_1_INVX1_211 gnd vdd FILL
XFILL_1_INVX1_222 gnd vdd FILL
XBUFX4_39 BUFX4_62/Y gnd DFFSR_84/R vdd BUFX4
XFILL_82_DFFSR_50 gnd vdd FILL
XFILL_82_DFFSR_61 gnd vdd FILL
XFILL_82_DFFSR_72 gnd vdd FILL
XFILL_82_DFFSR_83 gnd vdd FILL
XFILL_24_DFFSR_270 gnd vdd FILL
XFILL_82_DFFSR_94 gnd vdd FILL
XFILL_11_DFFSR_50 gnd vdd FILL
XFILL_5_INVX1_210 gnd vdd FILL
XFILL_21_MUX2X1_15 gnd vdd FILL
XFILL_11_DFFSR_61 gnd vdd FILL
XFILL_11_DFFSR_72 gnd vdd FILL
XFILL_21_MUX2X1_26 gnd vdd FILL
XFILL_5_INVX1_8 gnd vdd FILL
XFILL_21_MUX2X1_37 gnd vdd FILL
XFILL_5_INVX1_221 gnd vdd FILL
XFILL_11_DFFSR_83 gnd vdd FILL
XFILL_21_MUX2X1_48 gnd vdd FILL
XFILL_11_DFFSR_94 gnd vdd FILL
XFILL_21_MUX2X1_59 gnd vdd FILL
XFILL_16_7_2 gnd vdd FILL
XFILL_22_NOR3X1_2 gnd vdd FILL
XFILL_51_DFFSR_170 gnd vdd FILL
XFILL_15_2_1 gnd vdd FILL
XFILL_51_DFFSR_181 gnd vdd FILL
XFILL_51_DFFSR_60 gnd vdd FILL
XFILL_51_DFFSR_192 gnd vdd FILL
XFILL_51_DFFSR_71 gnd vdd FILL
XFILL_51_DFFSR_82 gnd vdd FILL
XFILL_51_DFFSR_93 gnd vdd FILL
XFILL_55_DFFSR_180 gnd vdd FILL
XFILL_55_DFFSR_191 gnd vdd FILL
XFILL_20_DFFSR_70 gnd vdd FILL
XFILL_9_MUX2X1_170 gnd vdd FILL
XFILL_20_DFFSR_81 gnd vdd FILL
XFILL_20_DFFSR_92 gnd vdd FILL
XFILL_5_NOR3X1_3 gnd vdd FILL
XFILL_9_MUX2X1_181 gnd vdd FILL
XFILL_59_DFFSR_190 gnd vdd FILL
XFILL_9_INVX8_2 gnd vdd FILL
XFILL_9_MUX2X1_192 gnd vdd FILL
XFILL_33_DFFSR_104 gnd vdd FILL
XFILL_33_DFFSR_115 gnd vdd FILL
XFILL_10_NAND2X1_6 gnd vdd FILL
XFILL_33_DFFSR_126 gnd vdd FILL
XFILL_33_DFFSR_137 gnd vdd FILL
XFILL_2_DFFSR_150 gnd vdd FILL
XFILL_2_DFFSR_161 gnd vdd FILL
XFILL_33_DFFSR_148 gnd vdd FILL
XFILL_60_DFFSR_80 gnd vdd FILL
XFILL_2_DFFSR_172 gnd vdd FILL
XFILL_33_DFFSR_159 gnd vdd FILL
XFILL_2_DFFSR_183 gnd vdd FILL
XFILL_60_DFFSR_91 gnd vdd FILL
XFILL_2_DFFSR_194 gnd vdd FILL
XFILL_37_DFFSR_103 gnd vdd FILL
XFILL_37_DFFSR_114 gnd vdd FILL
XFILL_37_DFFSR_125 gnd vdd FILL
XFILL_37_DFFSR_136 gnd vdd FILL
XFILL_11_NAND3X1_12 gnd vdd FILL
XFILL_37_DFFSR_147 gnd vdd FILL
XFILL_26_DFFSR_2 gnd vdd FILL
XFILL_6_DFFSR_160 gnd vdd FILL
XFILL_83_DFFSR_3 gnd vdd FILL
XFILL_37_DFFSR_158 gnd vdd FILL
XFILL_11_NAND3X1_23 gnd vdd FILL
XFILL_3_DFFSR_60 gnd vdd FILL
XFILL_6_DFFSR_171 gnd vdd FILL
XFILL_10_MUX2X1_80 gnd vdd FILL
XFILL_37_DFFSR_169 gnd vdd FILL
XFILL_11_NAND3X1_34 gnd vdd FILL
XFILL_3_DFFSR_71 gnd vdd FILL
XFILL_6_DFFSR_182 gnd vdd FILL
XFILL_3_DFFSR_82 gnd vdd FILL
XFILL_10_MUX2X1_91 gnd vdd FILL
XFILL_6_DFFSR_193 gnd vdd FILL
XFILL_11_NAND3X1_45 gnd vdd FILL
XFILL_3_DFFSR_93 gnd vdd FILL
XFILL_11_NAND3X1_56 gnd vdd FILL
XFILL_66_6_2 gnd vdd FILL
XFILL_31_CLKBUF1_12 gnd vdd FILL
XFILL_11_NAND3X1_67 gnd vdd FILL
XFILL_31_CLKBUF1_23 gnd vdd FILL
XFILL_11_NAND3X1_78 gnd vdd FILL
XFILL_31_CLKBUF1_34 gnd vdd FILL
XFILL_11_NAND3X1_89 gnd vdd FILL
XFILL_65_1_1 gnd vdd FILL
XFILL_14_MUX2X1_90 gnd vdd FILL
XFILL_2_NOR3X1_50 gnd vdd FILL
XFILL_83_DFFSR_204 gnd vdd FILL
XFILL_83_DFFSR_215 gnd vdd FILL
XFILL_10_DFFSR_8 gnd vdd FILL
XFILL_83_DFFSR_226 gnd vdd FILL
XFILL_83_DFFSR_237 gnd vdd FILL
XFILL_83_DFFSR_248 gnd vdd FILL
XFILL_83_DFFSR_259 gnd vdd FILL
XFILL_48_DFFSR_6 gnd vdd FILL
XFILL_87_DFFSR_203 gnd vdd FILL
XFILL_87_DFFSR_214 gnd vdd FILL
XFILL_87_DFFSR_225 gnd vdd FILL
XFILL_2_OAI22X1_19 gnd vdd FILL
XFILL_87_DFFSR_236 gnd vdd FILL
XFILL_87_DFFSR_247 gnd vdd FILL
XFILL_87_DFFSR_258 gnd vdd FILL
XFILL_22_DFFSR_180 gnd vdd FILL
XFILL_87_DFFSR_269 gnd vdd FILL
XFILL_22_DFFSR_191 gnd vdd FILL
XFILL_3_INVX1_120 gnd vdd FILL
XFILL_3_INVX1_131 gnd vdd FILL
XFILL_3_INVX1_142 gnd vdd FILL
XFILL_3_INVX1_153 gnd vdd FILL
XFILL_3_INVX1_164 gnd vdd FILL
XFILL_1_NAND3X1_40 gnd vdd FILL
XFILL_3_INVX1_175 gnd vdd FILL
XFILL_1_NAND3X1_51 gnd vdd FILL
XFILL_1_NAND3X1_62 gnd vdd FILL
XFILL_3_INVX1_186 gnd vdd FILL
XFILL_1_NAND3X1_73 gnd vdd FILL
XFILL_5_NAND2X1_20 gnd vdd FILL
XFILL_3_INVX1_197 gnd vdd FILL
XFILL_1_NAND3X1_84 gnd vdd FILL
XFILL_26_DFFSR_190 gnd vdd FILL
XFILL_5_NAND2X1_31 gnd vdd FILL
XFILL_5_NAND2X1_42 gnd vdd FILL
XFILL_1_NAND3X1_95 gnd vdd FILL
XFILL_5_NAND2X1_53 gnd vdd FILL
XFILL_7_INVX1_130 gnd vdd FILL
XFILL_7_INVX1_141 gnd vdd FILL
XFILL_5_NAND2X1_64 gnd vdd FILL
XFILL_7_INVX1_152 gnd vdd FILL
XFILL_5_NAND2X1_75 gnd vdd FILL
XFILL_5_NAND2X1_86 gnd vdd FILL
XFILL_7_INVX1_163 gnd vdd FILL
XFILL_7_INVX1_174 gnd vdd FILL
XFILL_7_INVX1_185 gnd vdd FILL
XFILL_7_INVX1_196 gnd vdd FILL
XFILL_13_CLKBUF1_17 gnd vdd FILL
XFILL_13_CLKBUF1_28 gnd vdd FILL
XFILL_13_CLKBUF1_39 gnd vdd FILL
XFILL_1_OAI22X1_4 gnd vdd FILL
XFILL_57_6_2 gnd vdd FILL
XFILL_56_1_1 gnd vdd FILL
XFILL_5_OAI22X1_3 gnd vdd FILL
XFILL_11_NOR2X1_102 gnd vdd FILL
XFILL_11_NOR2X1_113 gnd vdd FILL
XFILL_11_NOR2X1_124 gnd vdd FILL
XFILL_11_NOR2X1_135 gnd vdd FILL
XFILL_11_NOR2X1_146 gnd vdd FILL
XFILL_11_NOR2X1_157 gnd vdd FILL
XFILL_11_NOR2X1_168 gnd vdd FILL
XFILL_11_NOR2X1_179 gnd vdd FILL
XFILL_50_DFFSR_204 gnd vdd FILL
XFILL_50_DFFSR_215 gnd vdd FILL
XFILL_9_OAI22X1_2 gnd vdd FILL
XFILL_9_AOI21X1_20 gnd vdd FILL
XFILL_50_DFFSR_226 gnd vdd FILL
XFILL_50_DFFSR_237 gnd vdd FILL
XFILL_9_AOI21X1_31 gnd vdd FILL
XFILL_9_AOI21X1_42 gnd vdd FILL
XFILL_40_5_2 gnd vdd FILL
XFILL_50_DFFSR_248 gnd vdd FILL
XFILL_9_AOI21X1_53 gnd vdd FILL
XFILL_19_OAI22X1_11 gnd vdd FILL
XFILL_9_AOI21X1_64 gnd vdd FILL
XFILL_50_DFFSR_259 gnd vdd FILL
XFILL_19_OAI22X1_22 gnd vdd FILL
XFILL_9_AOI21X1_75 gnd vdd FILL
XFILL_19_OAI22X1_33 gnd vdd FILL
XFILL_19_OAI22X1_44 gnd vdd FILL
XFILL_54_DFFSR_203 gnd vdd FILL
XFILL_20_CLKBUF1_30 gnd vdd FILL
XFILL_20_CLKBUF1_41 gnd vdd FILL
XFILL_54_DFFSR_214 gnd vdd FILL
XFILL_54_DFFSR_225 gnd vdd FILL
XFILL_54_DFFSR_236 gnd vdd FILL
XFILL_54_DFFSR_247 gnd vdd FILL
XFILL_3_CLKBUF1_12 gnd vdd FILL
XFILL_54_DFFSR_258 gnd vdd FILL
XFILL_54_DFFSR_269 gnd vdd FILL
XFILL_3_CLKBUF1_23 gnd vdd FILL
XFILL_3_CLKBUF1_34 gnd vdd FILL
XFILL_58_DFFSR_202 gnd vdd FILL
XFILL_81_DFFSR_103 gnd vdd FILL
XFILL_58_DFFSR_213 gnd vdd FILL
XFILL_81_DFFSR_114 gnd vdd FILL
XFILL_11_MUX2X1_108 gnd vdd FILL
XFILL_11_MUX2X1_119 gnd vdd FILL
XFILL_81_DFFSR_125 gnd vdd FILL
XFILL_81_DFFSR_136 gnd vdd FILL
XFILL_58_DFFSR_224 gnd vdd FILL
XFILL_58_DFFSR_235 gnd vdd FILL
XFILL_58_DFFSR_246 gnd vdd FILL
XFILL_81_DFFSR_147 gnd vdd FILL
XFILL_6_BUFX2_1 gnd vdd FILL
XFILL_81_DFFSR_158 gnd vdd FILL
XFILL_58_DFFSR_257 gnd vdd FILL
XFILL_58_DFFSR_268 gnd vdd FILL
XFILL_81_DFFSR_169 gnd vdd FILL
XFILL_13_CLKBUF1_9 gnd vdd FILL
XFILL_1_DFFSR_206 gnd vdd FILL
XFILL_85_DFFSR_102 gnd vdd FILL
XFILL_74_DFFSR_19 gnd vdd FILL
XFILL_12_OAI21X1_13 gnd vdd FILL
XFILL_1_DFFSR_217 gnd vdd FILL
XFILL_85_DFFSR_113 gnd vdd FILL
XFILL_85_DFFSR_124 gnd vdd FILL
XFILL_12_OAI21X1_24 gnd vdd FILL
XFILL_1_DFFSR_228 gnd vdd FILL
XFILL_85_DFFSR_135 gnd vdd FILL
XFILL_1_DFFSR_239 gnd vdd FILL
XFILL_1_NOR2X1_130 gnd vdd FILL
XFILL_85_DFFSR_146 gnd vdd FILL
XFILL_1_NOR2X1_141 gnd vdd FILL
XFILL_12_OAI21X1_35 gnd vdd FILL
XFILL_12_OAI21X1_46 gnd vdd FILL
XFILL_1_NOR2X1_152 gnd vdd FILL
XFILL_17_MUX2X1_9 gnd vdd FILL
XFILL_85_DFFSR_157 gnd vdd FILL
XFILL_85_DFFSR_168 gnd vdd FILL
XFILL_1_NOR2X1_163 gnd vdd FILL
XFILL_85_DFFSR_179 gnd vdd FILL
XFILL_17_CLKBUF1_8 gnd vdd FILL
XFILL_1_NOR2X1_174 gnd vdd FILL
XFILL_5_DFFSR_205 gnd vdd FILL
XFILL_1_NOR2X1_185 gnd vdd FILL
XFILL_2_NAND3X1_5 gnd vdd FILL
XFILL_1_NOR2X1_196 gnd vdd FILL
XFILL_8_BUFX4_20 gnd vdd FILL
XFILL_48_6_2 gnd vdd FILL
XFILL_5_DFFSR_216 gnd vdd FILL
XFILL_8_BUFX4_31 gnd vdd FILL
XFILL_5_DFFSR_227 gnd vdd FILL
XFILL_8_BUFX4_42 gnd vdd FILL
XFILL_5_DFFSR_238 gnd vdd FILL
XFILL_47_1_1 gnd vdd FILL
XFILL_8_BUFX4_53 gnd vdd FILL
XFILL_5_DFFSR_249 gnd vdd FILL
XFILL_8_BUFX4_64 gnd vdd FILL
XFILL_43_DFFSR_18 gnd vdd FILL
XFILL_13_BUFX4_103 gnd vdd FILL
XFILL_43_DFFSR_29 gnd vdd FILL
XFILL_8_BUFX4_75 gnd vdd FILL
XFILL_8_BUFX4_86 gnd vdd FILL
XFILL_8_BUFX4_97 gnd vdd FILL
XFILL_9_OAI22X1_50 gnd vdd FILL
XFILL_9_DFFSR_204 gnd vdd FILL
XFILL_9_DFFSR_215 gnd vdd FILL
XFILL_6_NAND3X1_4 gnd vdd FILL
XFILL_9_DFFSR_226 gnd vdd FILL
XFILL_9_DFFSR_237 gnd vdd FILL
XFILL_9_DFFSR_248 gnd vdd FILL
XFILL_9_DFFSR_259 gnd vdd FILL
XFILL_83_DFFSR_17 gnd vdd FILL
XFILL_83_DFFSR_28 gnd vdd FILL
XFILL_1_MUX2X1_103 gnd vdd FILL
XFILL_83_DFFSR_39 gnd vdd FILL
XFILL_1_MUX2X1_114 gnd vdd FILL
XFILL_1_MUX2X1_125 gnd vdd FILL
XFILL_12_DFFSR_17 gnd vdd FILL
XNAND3X1_130 DFFSR_159/Q BUFX4_88/Y NOR2X1_36/Y gnd OAI21X1_22/C vdd NAND3X1
XFILL_31_5_2 gnd vdd FILL
XFILL_12_DFFSR_28 gnd vdd FILL
XFILL_1_MUX2X1_136 gnd vdd FILL
XFILL_12_DFFSR_39 gnd vdd FILL
XFILL_1_MUX2X1_147 gnd vdd FILL
XFILL_1_MUX2X1_158 gnd vdd FILL
XFILL_30_0_1 gnd vdd FILL
XFILL_87_DFFSR_4 gnd vdd FILL
XFILL_1_MUX2X1_169 gnd vdd FILL
XFILL_6_INVX2_1 gnd vdd FILL
XFILL_70_DFFSR_190 gnd vdd FILL
XFILL_52_DFFSR_16 gnd vdd FILL
XFILL_2_OAI21X1_30 gnd vdd FILL
XFILL_21_DFFSR_203 gnd vdd FILL
XFILL_52_DFFSR_27 gnd vdd FILL
XFILL_2_OAI21X1_41 gnd vdd FILL
XFILL_52_DFFSR_38 gnd vdd FILL
XFILL_21_DFFSR_214 gnd vdd FILL
XFILL_11_NOR2X1_16 gnd vdd FILL
XFILL_11_NOR2X1_27 gnd vdd FILL
XFILL_52_DFFSR_49 gnd vdd FILL
XFILL_21_DFFSR_225 gnd vdd FILL
XFILL_21_DFFSR_236 gnd vdd FILL
XFILL_11_NOR2X1_38 gnd vdd FILL
XFILL_21_DFFSR_247 gnd vdd FILL
XFILL_21_DFFSR_258 gnd vdd FILL
XFILL_11_NOR2X1_49 gnd vdd FILL
XFILL_21_DFFSR_269 gnd vdd FILL
XFILL_25_DFFSR_202 gnd vdd FILL
XFILL_2_INVX1_209 gnd vdd FILL
XFILL_25_DFFSR_213 gnd vdd FILL
XFILL_9_MUX2X1_8 gnd vdd FILL
XFILL_6_AOI22X1_9 gnd vdd FILL
XFILL_25_DFFSR_224 gnd vdd FILL
XFILL_14_DFFSR_9 gnd vdd FILL
XFILL_25_DFFSR_235 gnd vdd FILL
XFILL_21_DFFSR_15 gnd vdd FILL
XFILL_21_DFFSR_26 gnd vdd FILL
XFILL_25_DFFSR_246 gnd vdd FILL
XFILL_25_DFFSR_257 gnd vdd FILL
XFILL_21_DFFSR_37 gnd vdd FILL
XFILL_25_DFFSR_268 gnd vdd FILL
XFILL_21_DFFSR_48 gnd vdd FILL
XFILL_6_INVX1_208 gnd vdd FILL
XFILL_12_BUFX4_80 gnd vdd FILL
XFILL_21_DFFSR_59 gnd vdd FILL
XFILL_29_DFFSR_201 gnd vdd FILL
XFILL_52_DFFSR_102 gnd vdd FILL
XFILL_12_BUFX4_91 gnd vdd FILL
XFILL_29_DFFSR_212 gnd vdd FILL
XFILL_6_INVX1_219 gnd vdd FILL
XFILL_52_DFFSR_113 gnd vdd FILL
XFILL_52_DFFSR_124 gnd vdd FILL
XFILL_52_DFFSR_135 gnd vdd FILL
XFILL_29_DFFSR_223 gnd vdd FILL
XFILL_29_DFFSR_234 gnd vdd FILL
XFILL_61_DFFSR_14 gnd vdd FILL
XFILL_52_DFFSR_146 gnd vdd FILL
XFILL_61_DFFSR_25 gnd vdd FILL
XFILL_29_DFFSR_245 gnd vdd FILL
XFILL_52_DFFSR_157 gnd vdd FILL
XFILL_39_6_2 gnd vdd FILL
XFILL_61_DFFSR_36 gnd vdd FILL
XFILL_29_DFFSR_256 gnd vdd FILL
XFILL_29_DFFSR_267 gnd vdd FILL
XFILL_52_DFFSR_168 gnd vdd FILL
XFILL_52_DFFSR_179 gnd vdd FILL
XFILL_61_DFFSR_47 gnd vdd FILL
XFILL_56_DFFSR_101 gnd vdd FILL
XFILL_61_DFFSR_58 gnd vdd FILL
XFILL_38_1_1 gnd vdd FILL
XFILL_61_DFFSR_69 gnd vdd FILL
XFILL_56_DFFSR_112 gnd vdd FILL
XFILL_4_NAND3X1_17 gnd vdd FILL
XFILL_56_DFFSR_123 gnd vdd FILL
XFILL_56_DFFSR_134 gnd vdd FILL
XFILL_4_NAND3X1_28 gnd vdd FILL
XFILL_56_DFFSR_145 gnd vdd FILL
XFILL_4_NAND3X1_39 gnd vdd FILL
XFILL_56_DFFSR_156 gnd vdd FILL
XFILL_4_DFFSR_16 gnd vdd FILL
XFILL_56_DFFSR_167 gnd vdd FILL
XFILL_4_DFFSR_27 gnd vdd FILL
XFILL_56_DFFSR_178 gnd vdd FILL
XFILL_8_NAND2X1_19 gnd vdd FILL
XFILL_30_DFFSR_13 gnd vdd FILL
XFILL_4_DFFSR_38 gnd vdd FILL
XFILL_56_DFFSR_189 gnd vdd FILL
XFILL_30_DFFSR_24 gnd vdd FILL
XFILL_4_DFFSR_49 gnd vdd FILL
XFILL_30_DFFSR_35 gnd vdd FILL
XFILL_30_DFFSR_46 gnd vdd FILL
XFILL_30_DFFSR_57 gnd vdd FILL
XFILL_30_DFFSR_68 gnd vdd FILL
XFILL_30_DFFSR_79 gnd vdd FILL
XFILL_6_INVX1_70 gnd vdd FILL
XFILL_18_MUX2X1_150 gnd vdd FILL
XFILL_22_5_2 gnd vdd FILL
XFILL_6_INVX1_81 gnd vdd FILL
XFILL_6_INVX1_92 gnd vdd FILL
XFILL_18_MUX2X1_161 gnd vdd FILL
XFILL_3_DFFSR_104 gnd vdd FILL
XFILL_70_DFFSR_12 gnd vdd FILL
XFILL_21_0_1 gnd vdd FILL
XFILL_3_DFFSR_115 gnd vdd FILL
XFILL_18_MUX2X1_172 gnd vdd FILL
XFILL_70_DFFSR_23 gnd vdd FILL
XFILL_3_DFFSR_126 gnd vdd FILL
XFILL_70_DFFSR_34 gnd vdd FILL
XFILL_18_MUX2X1_183 gnd vdd FILL
XFILL_3_DFFSR_137 gnd vdd FILL
XFILL_18_MUX2X1_194 gnd vdd FILL
XFILL_70_DFFSR_45 gnd vdd FILL
XFILL_70_DFFSR_56 gnd vdd FILL
XFILL_13_MUX2X1_2 gnd vdd FILL
XFILL_3_DFFSR_148 gnd vdd FILL
XFILL_70_DFFSR_67 gnd vdd FILL
XFILL_3_DFFSR_159 gnd vdd FILL
XFILL_70_DFFSR_78 gnd vdd FILL
XFILL_70_DFFSR_89 gnd vdd FILL
XFILL_7_DFFSR_103 gnd vdd FILL
XFILL_7_DFFSR_114 gnd vdd FILL
XFILL_11_MUX2X1_12 gnd vdd FILL
XFILL_11_MUX2X1_23 gnd vdd FILL
XFILL_7_DFFSR_125 gnd vdd FILL
XFILL_7_DFFSR_136 gnd vdd FILL
XDFFSR_150 DFFSR_150/Q DFFSR_58/CLK DFFSR_91/R vdd DFFSR_150/D gnd vdd DFFSR
XFILL_11_MUX2X1_34 gnd vdd FILL
XDFFSR_161 INVX1_146/A DFFSR_70/CLK DFFSR_98/R vdd MUX2X1_79/Y gnd vdd DFFSR
XFILL_11_MUX2X1_45 gnd vdd FILL
XFILL_7_DFFSR_147 gnd vdd FILL
XBUFX4_2 BUFX4_2/A gnd BUFX4_2/Y vdd BUFX4
XFILL_7_DFFSR_158 gnd vdd FILL
XDFFSR_172 NOR2X1_2/A DFFSR_58/CLK DFFSR_23/R vdd DFFSR_172/D gnd vdd DFFSR
XFILL_11_MUX2X1_56 gnd vdd FILL
XDFFSR_183 INVX1_143/A DFFSR_99/CLK DFFSR_99/R vdd DFFSR_183/D gnd vdd DFFSR
XFILL_7_DFFSR_169 gnd vdd FILL
XFILL_11_MUX2X1_67 gnd vdd FILL
XFILL_10_NOR3X1_8 gnd vdd FILL
XFILL_11_MUX2X1_78 gnd vdd FILL
XFILL_4_BUFX4_90 gnd vdd FILL
XDFFSR_194 INVX1_130/A DFFSR_1/CLK DFFSR_1/R vdd DFFSR_194/D gnd vdd DFFSR
XFILL_11_MUX2X1_89 gnd vdd FILL
XFILL_15_MUX2X1_11 gnd vdd FILL
XFILL_15_MUX2X1_22 gnd vdd FILL
XFILL_15_MUX2X1_33 gnd vdd FILL
XFILL_15_MUX2X1_44 gnd vdd FILL
XFILL_15_MUX2X1_55 gnd vdd FILL
XFILL_15_MUX2X1_66 gnd vdd FILL
XFILL_15_MUX2X1_77 gnd vdd FILL
XFILL_3_NOR3X1_15 gnd vdd FILL
XFILL_15_MUX2X1_88 gnd vdd FILL
XFILL_15_MUX2X1_99 gnd vdd FILL
XFILL_3_NOR3X1_26 gnd vdd FILL
XFILL_19_MUX2X1_10 gnd vdd FILL
XFILL_3_NOR3X1_37 gnd vdd FILL
XFILL_19_MUX2X1_21 gnd vdd FILL
XFILL_3_NOR3X1_48 gnd vdd FILL
XFILL_23_CLKBUF1_18 gnd vdd FILL
XFILL_19_MUX2X1_32 gnd vdd FILL
XFILL_23_CLKBUF1_29 gnd vdd FILL
XFILL_5_6_2 gnd vdd FILL
XFILL_19_MUX2X1_43 gnd vdd FILL
XFILL_19_MUX2X1_54 gnd vdd FILL
XFILL_6_NOR2X1_3 gnd vdd FILL
XFILL_29_1_1 gnd vdd FILL
XFILL_4_1_1 gnd vdd FILL
XFILL_19_MUX2X1_65 gnd vdd FILL
XFILL_7_NOR3X1_14 gnd vdd FILL
XFILL_19_MUX2X1_76 gnd vdd FILL
XFILL_19_MUX2X1_87 gnd vdd FILL
XFILL_7_NOR3X1_25 gnd vdd FILL
XFILL_19_MUX2X1_98 gnd vdd FILL
XNOR3X1_50 NOR3X1_50/A NOR3X1_50/B NOR3X1_50/C gnd NOR3X1_50/Y vdd NOR3X1
XFILL_0_INVX1_108 gnd vdd FILL
XFILL_7_NOR3X1_36 gnd vdd FILL
XFILL_23_DFFSR_101 gnd vdd FILL
XFILL_7_NOR3X1_47 gnd vdd FILL
XFILL_0_INVX1_119 gnd vdd FILL
XFILL_23_DFFSR_112 gnd vdd FILL
XFILL_23_DFFSR_123 gnd vdd FILL
XFILL_23_DFFSR_134 gnd vdd FILL
XFILL_1_AOI21X1_19 gnd vdd FILL
XFILL_23_DFFSR_145 gnd vdd FILL
XFILL_23_DFFSR_156 gnd vdd FILL
XFILL_23_DFFSR_167 gnd vdd FILL
XFILL_23_DFFSR_178 gnd vdd FILL
XFILL_5_MUX2X1_1 gnd vdd FILL
XFILL_4_INVX1_107 gnd vdd FILL
XFILL_27_DFFSR_100 gnd vdd FILL
XFILL_23_DFFSR_189 gnd vdd FILL
XFILL_4_INVX1_118 gnd vdd FILL
XFILL_4_INVX1_129 gnd vdd FILL
XFILL_27_DFFSR_111 gnd vdd FILL
XFILL_4_NOR2X1_107 gnd vdd FILL
XFILL_13_5_2 gnd vdd FILL
XFILL_27_DFFSR_122 gnd vdd FILL
XFILL_31_DFFSR_3 gnd vdd FILL
XFILL_4_NOR2X1_118 gnd vdd FILL
XFILL_27_DFFSR_133 gnd vdd FILL
XFILL_27_DFFSR_144 gnd vdd FILL
XFILL_4_NOR2X1_129 gnd vdd FILL
XFILL_10_NAND3X1_20 gnd vdd FILL
XFILL_27_DFFSR_155 gnd vdd FILL
XFILL_12_0_1 gnd vdd FILL
XFILL_10_NAND3X1_31 gnd vdd FILL
XFILL_27_DFFSR_166 gnd vdd FILL
XFILL_27_DFFSR_177 gnd vdd FILL
XFILL_10_NAND3X1_42 gnd vdd FILL
XFILL_10_NAND3X1_53 gnd vdd FILL
XFILL_27_DFFSR_188 gnd vdd FILL
XFILL_69_DFFSR_1 gnd vdd FILL
XFILL_10_NAND3X1_64 gnd vdd FILL
XFILL_27_DFFSR_199 gnd vdd FILL
XFILL_30_CLKBUF1_20 gnd vdd FILL
XFILL_10_NAND3X1_75 gnd vdd FILL
XFILL_2_NOR3X1_7 gnd vdd FILL
XFILL_10_NAND3X1_86 gnd vdd FILL
XFILL_30_CLKBUF1_31 gnd vdd FILL
XFILL_10_NAND3X1_97 gnd vdd FILL
XFILL_30_CLKBUF1_42 gnd vdd FILL
XFILL_23_NOR3X1_12 gnd vdd FILL
XFILL_39_DFFSR_90 gnd vdd FILL
XFILL_23_NOR3X1_23 gnd vdd FILL
XFILL_23_NOR3X1_34 gnd vdd FILL
XFILL_73_DFFSR_201 gnd vdd FILL
XFILL_23_NOR3X1_45 gnd vdd FILL
XFILL_21_MUX2X1_109 gnd vdd FILL
XFILL_73_DFFSR_212 gnd vdd FILL
XFILL_73_DFFSR_223 gnd vdd FILL
XFILL_0_DFFSR_20 gnd vdd FILL
XFILL_73_DFFSR_234 gnd vdd FILL
XFILL_0_DFFSR_31 gnd vdd FILL
XFILL_0_DFFSR_42 gnd vdd FILL
XFILL_73_DFFSR_245 gnd vdd FILL
XFILL_27_NOR3X1_11 gnd vdd FILL
XFILL_73_DFFSR_256 gnd vdd FILL
XFILL_73_DFFSR_267 gnd vdd FILL
XFILL_0_DFFSR_53 gnd vdd FILL
XFILL_27_NOR3X1_22 gnd vdd FILL
XFILL_27_NOR3X1_33 gnd vdd FILL
XFILL_0_DFFSR_64 gnd vdd FILL
XFILL_53_DFFSR_7 gnd vdd FILL
XFILL_0_DFFSR_75 gnd vdd FILL
XFILL_0_DFFSR_86 gnd vdd FILL
XFILL_77_DFFSR_200 gnd vdd FILL
XFILL_27_NOR3X1_44 gnd vdd FILL
XFILL_7_5 gnd vdd FILL
XFILL_77_DFFSR_211 gnd vdd FILL
XFILL_0_DFFSR_97 gnd vdd FILL
XFILL_77_DFFSR_222 gnd vdd FILL
XFILL_1_OAI22X1_16 gnd vdd FILL
XFILL_77_DFFSR_233 gnd vdd FILL
XFILL_77_DFFSR_244 gnd vdd FILL
XFILL_1_OAI22X1_27 gnd vdd FILL
XFILL_63_7 gnd vdd FILL
XFILL_77_DFFSR_255 gnd vdd FILL
XFILL_1_OAI22X1_38 gnd vdd FILL
XFILL_77_DFFSR_266 gnd vdd FILL
XFILL_1_OAI22X1_49 gnd vdd FILL
XFILL_32_CLKBUF1_7 gnd vdd FILL
XFILL_5_OAI21X1_18 gnd vdd FILL
XFILL_5_OAI21X1_29 gnd vdd FILL
XFILL_63_4_2 gnd vdd FILL
XFILL_0_NAND3X1_70 gnd vdd FILL
XFILL_0_NAND3X1_81 gnd vdd FILL
XFILL_0_NAND3X1_92 gnd vdd FILL
XFILL_4_NAND2X1_50 gnd vdd FILL
XFILL_4_NAND2X1_61 gnd vdd FILL
XFILL_4_NAND2X1_72 gnd vdd FILL
XFILL_4_NAND2X1_83 gnd vdd FILL
XFILL_4_NAND2X1_94 gnd vdd FILL
XFILL_12_CLKBUF1_14 gnd vdd FILL
XFILL_12_CLKBUF1_25 gnd vdd FILL
XFILL_12_CLKBUF1_36 gnd vdd FILL
XFILL_10_NOR2X1_110 gnd vdd FILL
XFILL_10_NOR2X1_121 gnd vdd FILL
XFILL_10_NOR2X1_132 gnd vdd FILL
XFILL_10_NOR2X1_143 gnd vdd FILL
XFILL_10_NOR2X1_154 gnd vdd FILL
XFILL_10_NOR2X1_165 gnd vdd FILL
XFILL_40_DFFSR_201 gnd vdd FILL
XFILL_10_NOR2X1_176 gnd vdd FILL
XFILL_10_NOR2X1_187 gnd vdd FILL
XFILL_2_OAI21X1_2 gnd vdd FILL
XFILL_40_DFFSR_212 gnd vdd FILL
XFILL_10_NOR2X1_198 gnd vdd FILL
XFILL_40_DFFSR_223 gnd vdd FILL
XFILL_40_DFFSR_234 gnd vdd FILL
XFILL_40_DFFSR_245 gnd vdd FILL
XFILL_8_AOI21X1_50 gnd vdd FILL
XFILL_40_DFFSR_256 gnd vdd FILL
XNAND3X1_5 DFFSR_18/Q BUFX4_8/Y NOR2X1_36/Y gnd NAND3X1_8/B vdd NAND3X1
XFILL_8_AOI21X1_61 gnd vdd FILL
XFILL_40_DFFSR_267 gnd vdd FILL
XFILL_8_AOI21X1_72 gnd vdd FILL
XFILL_18_OAI22X1_30 gnd vdd FILL
XFILL_18_OAI22X1_41 gnd vdd FILL
XFILL_44_DFFSR_200 gnd vdd FILL
XFILL_44_DFFSR_211 gnd vdd FILL
XFILL_6_OAI21X1_1 gnd vdd FILL
XFILL_44_DFFSR_222 gnd vdd FILL
XFILL_44_DFFSR_233 gnd vdd FILL
XFILL_44_DFFSR_244 gnd vdd FILL
XFILL_44_DFFSR_255 gnd vdd FILL
XFILL_2_CLKBUF1_20 gnd vdd FILL
XFILL_3_NOR2X1_70 gnd vdd FILL
XFILL_44_DFFSR_266 gnd vdd FILL
XFILL_13_BUFX4_14 gnd vdd FILL
XFILL_3_NOR2X1_81 gnd vdd FILL
XFILL_13_BUFX4_25 gnd vdd FILL
XFILL_3_NOR2X1_92 gnd vdd FILL
XFILL_2_CLKBUF1_31 gnd vdd FILL
XFILL_13_BUFX4_36 gnd vdd FILL
XFILL_13_BUFX4_47 gnd vdd FILL
XFILL_71_DFFSR_100 gnd vdd FILL
XFILL_2_CLKBUF1_42 gnd vdd FILL
XFILL_54_4_2 gnd vdd FILL
XFILL_48_DFFSR_210 gnd vdd FILL
XFILL_71_DFFSR_111 gnd vdd FILL
XFILL_10_MUX2X1_105 gnd vdd FILL
XFILL_10_MUX2X1_116 gnd vdd FILL
XFILL_48_DFFSR_221 gnd vdd FILL
XFILL_71_DFFSR_122 gnd vdd FILL
XFILL_13_BUFX4_58 gnd vdd FILL
XFILL_71_DFFSR_133 gnd vdd FILL
XFILL_13_BUFX4_69 gnd vdd FILL
XFILL_10_MUX2X1_127 gnd vdd FILL
XFILL_71_DFFSR_144 gnd vdd FILL
XFILL_10_MUX2X1_138 gnd vdd FILL
XFILL_48_DFFSR_232 gnd vdd FILL
XFILL_48_DFFSR_243 gnd vdd FILL
XFILL_10_MUX2X1_149 gnd vdd FILL
XFILL_71_DFFSR_155 gnd vdd FILL
XFILL_48_DFFSR_254 gnd vdd FILL
XFILL_71_DFFSR_166 gnd vdd FILL
XFILL_48_DFFSR_265 gnd vdd FILL
XFILL_71_DFFSR_177 gnd vdd FILL
XFILL_7_NOR2X1_80 gnd vdd FILL
XFILL_71_DFFSR_188 gnd vdd FILL
XFILL_7_NOR2X1_91 gnd vdd FILL
XFILL_71_DFFSR_199 gnd vdd FILL
XFILL_11_OAI21X1_10 gnd vdd FILL
XFILL_75_DFFSR_110 gnd vdd FILL
XFILL_11_OAI21X1_21 gnd vdd FILL
XFILL_75_DFFSR_121 gnd vdd FILL
XFILL_75_DFFSR_132 gnd vdd FILL
XFILL_11_OAI21X1_32 gnd vdd FILL
XFILL_0_DFFSR_2 gnd vdd FILL
XFILL_75_DFFSR_143 gnd vdd FILL
XFILL_75_DFFSR_154 gnd vdd FILL
XFILL_11_OAI21X1_43 gnd vdd FILL
XFILL_0_NOR2X1_160 gnd vdd FILL
XFILL_75_DFFSR_165 gnd vdd FILL
XFILL_0_NOR2X1_171 gnd vdd FILL
XFILL_70_DFFSR_1 gnd vdd FILL
XFILL_75_DFFSR_176 gnd vdd FILL
XFILL_75_DFFSR_187 gnd vdd FILL
XFILL_0_NOR2X1_182 gnd vdd FILL
XFILL_75_DFFSR_198 gnd vdd FILL
XFILL_0_NOR2X1_193 gnd vdd FILL
XFILL_79_DFFSR_120 gnd vdd FILL
XFILL_79_DFFSR_131 gnd vdd FILL
XFILL_79_DFFSR_142 gnd vdd FILL
XFILL_79_DFFSR_153 gnd vdd FILL
XFILL_7_INVX1_15 gnd vdd FILL
XFILL_7_INVX1_26 gnd vdd FILL
XFILL_79_DFFSR_164 gnd vdd FILL
XFILL_7_INVX1_37 gnd vdd FILL
XFILL_79_DFFSR_175 gnd vdd FILL
XINVX1_209 DFFSR_78/Q gnd INVX1_209/Y vdd INVX1
XFILL_79_DFFSR_186 gnd vdd FILL
XFILL_7_INVX1_48 gnd vdd FILL
XFILL_8_AND2X2_7 gnd vdd FILL
XFILL_79_DFFSR_197 gnd vdd FILL
XFILL_7_INVX1_59 gnd vdd FILL
XFILL_0_MUX2X1_100 gnd vdd FILL
XFILL_0_MUX2X1_111 gnd vdd FILL
XFILL_0_MUX2X1_122 gnd vdd FILL
XFILL_3_NAND2X1_3 gnd vdd FILL
XFILL_35_DFFSR_4 gnd vdd FILL
XFILL_0_MUX2X1_133 gnd vdd FILL
XFILL_5_BUFX4_13 gnd vdd FILL
XFILL_0_MUX2X1_144 gnd vdd FILL
XFILL_0_MUX2X1_155 gnd vdd FILL
XFILL_13_NAND3X1_19 gnd vdd FILL
XFILL_5_BUFX4_24 gnd vdd FILL
XFILL_0_MUX2X1_166 gnd vdd FILL
XFILL_5_BUFX4_35 gnd vdd FILL
XFILL_5_BUFX4_46 gnd vdd FILL
XFILL_0_MUX2X1_177 gnd vdd FILL
XFILL_5_BUFX4_57 gnd vdd FILL
XFILL_0_MUX2X1_188 gnd vdd FILL
XFILL_5_BUFX4_68 gnd vdd FILL
XFILL_7_NAND2X1_2 gnd vdd FILL
XFILL_11_DFFSR_200 gnd vdd FILL
XFILL_5_BUFX4_79 gnd vdd FILL
XFILL_33_CLKBUF1_19 gnd vdd FILL
XFILL_11_DFFSR_211 gnd vdd FILL
XFILL_11_DFFSR_222 gnd vdd FILL
XFILL_11_DFFSR_233 gnd vdd FILL
XFILL_11_DFFSR_244 gnd vdd FILL
XFILL_11_DFFSR_255 gnd vdd FILL
XFILL_45_4_2 gnd vdd FILL
XFILL_11_DFFSR_266 gnd vdd FILL
XFILL_15_DFFSR_210 gnd vdd FILL
XFILL_15_DFFSR_221 gnd vdd FILL
XFILL_15_DFFSR_232 gnd vdd FILL
XFILL_15_DFFSR_243 gnd vdd FILL
XFILL_15_DFFSR_254 gnd vdd FILL
XFILL_15_DFFSR_265 gnd vdd FILL
XFILL_57_DFFSR_8 gnd vdd FILL
XFILL_12_AND2X2_1 gnd vdd FILL
XFILL_42_DFFSR_110 gnd vdd FILL
XFILL_19_DFFSR_220 gnd vdd FILL
XFILL_42_DFFSR_121 gnd vdd FILL
XFILL_42_DFFSR_132 gnd vdd FILL
XFILL_3_AOI21X1_8 gnd vdd FILL
XFILL_42_DFFSR_143 gnd vdd FILL
XFILL_19_DFFSR_231 gnd vdd FILL
XFILL_19_DFFSR_242 gnd vdd FILL
XFILL_42_DFFSR_154 gnd vdd FILL
XFILL_19_DFFSR_253 gnd vdd FILL
XFILL_42_DFFSR_165 gnd vdd FILL
XFILL_19_DFFSR_264 gnd vdd FILL
XFILL_19_DFFSR_275 gnd vdd FILL
XFILL_42_DFFSR_176 gnd vdd FILL
XFILL_42_DFFSR_187 gnd vdd FILL
XFILL_42_DFFSR_198 gnd vdd FILL
XFILL_46_DFFSR_120 gnd vdd FILL
XFILL_3_NAND3X1_14 gnd vdd FILL
XFILL_46_DFFSR_131 gnd vdd FILL
XFILL_7_AOI21X1_7 gnd vdd FILL
XFILL_3_NAND3X1_25 gnd vdd FILL
XFILL_46_DFFSR_142 gnd vdd FILL
XFILL_3_NAND3X1_36 gnd vdd FILL
XFILL_46_DFFSR_153 gnd vdd FILL
XNOR3X1_8 NOR3X1_8/A NOR3X1_8/B NOR3X1_8/C gnd NOR3X1_8/Y vdd NOR3X1
XFILL_3_NAND3X1_47 gnd vdd FILL
XFILL_3_NAND3X1_58 gnd vdd FILL
XFILL_7_NAND2X1_16 gnd vdd FILL
XFILL_46_DFFSR_164 gnd vdd FILL
XFILL_3_NAND3X1_69 gnd vdd FILL
XFILL_46_DFFSR_175 gnd vdd FILL
XFILL_7_NAND2X1_27 gnd vdd FILL
XFILL_46_DFFSR_186 gnd vdd FILL
XFILL_46_DFFSR_197 gnd vdd FILL
XFILL_7_NAND2X1_38 gnd vdd FILL
XFILL_7_NAND2X1_49 gnd vdd FILL
XFILL_12_AOI22X1_4 gnd vdd FILL
XMUX2X1_190 BUFX4_72/Y INVX1_10/Y NOR2X1_169/Y gnd DFFSR_52/D vdd MUX2X1
XFILL_5_2 gnd vdd FILL
XFILL_17_MUX2X1_180 gnd vdd FILL
XFILL_17_MUX2X1_191 gnd vdd FILL
XFILL_61_4 gnd vdd FILL
XFILL_16_AOI22X1_3 gnd vdd FILL
XFILL_54_3 gnd vdd FILL
XFILL_28_DFFSR_109 gnd vdd FILL
XFILL_64_7_0 gnd vdd FILL
XFILL_11_NOR2X1_8 gnd vdd FILL
XFILL_36_4_2 gnd vdd FILL
XFILL_3_INVX1_30 gnd vdd FILL
XFILL_3_INVX1_41 gnd vdd FILL
XFILL_3_INVX1_52 gnd vdd FILL
XFILL_3_INVX1_63 gnd vdd FILL
XFILL_49_DFFSR_11 gnd vdd FILL
XFILL_3_INVX1_74 gnd vdd FILL
XFILL_3_INVX1_85 gnd vdd FILL
XFILL_3_INVX1_96 gnd vdd FILL
XFILL_49_DFFSR_22 gnd vdd FILL
XFILL_49_DFFSR_33 gnd vdd FILL
XFILL_49_DFFSR_44 gnd vdd FILL
XFILL_49_DFFSR_55 gnd vdd FILL
XFILL_49_DFFSR_66 gnd vdd FILL
XFILL_10_MUX2X1_6 gnd vdd FILL
XFILL_49_DFFSR_77 gnd vdd FILL
XFILL_49_DFFSR_88 gnd vdd FILL
XFILL_49_DFFSR_99 gnd vdd FILL
XFILL_22_CLKBUF1_15 gnd vdd FILL
XFILL_22_CLKBUF1_26 gnd vdd FILL
XFILL_22_CLKBUF1_37 gnd vdd FILL
XFILL_18_DFFSR_10 gnd vdd FILL
XFILL_18_DFFSR_21 gnd vdd FILL
XFILL_1_BUFX4_50 gnd vdd FILL
XFILL_1_BUFX4_61 gnd vdd FILL
XFILL_1_BUFX4_72 gnd vdd FILL
XFILL_18_DFFSR_32 gnd vdd FILL
XFILL_5_CLKBUF1_19 gnd vdd FILL
XFILL_1_BUFX4_83 gnd vdd FILL
XFILL_18_DFFSR_43 gnd vdd FILL
XFILL_18_DFFSR_54 gnd vdd FILL
XFILL_18_DFFSR_65 gnd vdd FILL
XFILL_1_BUFX4_94 gnd vdd FILL
XFILL_18_DFFSR_76 gnd vdd FILL
XFILL_0_AOI21X1_16 gnd vdd FILL
XFILL_13_DFFSR_120 gnd vdd FILL
XFILL_78_DFFSR_209 gnd vdd FILL
XFILL_13_DFFSR_131 gnd vdd FILL
XFILL_18_DFFSR_87 gnd vdd FILL
XFILL_18_DFFSR_98 gnd vdd FILL
XFILL_13_DFFSR_142 gnd vdd FILL
XFILL_0_AOI21X1_27 gnd vdd FILL
XFILL_13_DFFSR_153 gnd vdd FILL
XFILL_58_DFFSR_20 gnd vdd FILL
XFILL_0_AOI21X1_38 gnd vdd FILL
XFILL_0_AOI21X1_49 gnd vdd FILL
XFILL_58_DFFSR_31 gnd vdd FILL
XFILL_29_NOR3X1_6 gnd vdd FILL
XFILL_13_DFFSR_164 gnd vdd FILL
XFILL_2_CLKBUF1_7 gnd vdd FILL
XFILL_13_DFFSR_175 gnd vdd FILL
XFILL_10_OAI22X1_18 gnd vdd FILL
XFILL_58_DFFSR_42 gnd vdd FILL
XFILL_13_DFFSR_186 gnd vdd FILL
XFILL_10_OAI22X1_29 gnd vdd FILL
XFILL_58_DFFSR_53 gnd vdd FILL
XFILL_13_DFFSR_197 gnd vdd FILL
XFILL_58_DFFSR_64 gnd vdd FILL
XFILL_3_NOR2X1_104 gnd vdd FILL
XFILL_58_DFFSR_75 gnd vdd FILL
XFILL_58_DFFSR_86 gnd vdd FILL
XFILL_17_DFFSR_130 gnd vdd FILL
XFILL_3_NOR2X1_115 gnd vdd FILL
XFILL_4_DFFSR_3 gnd vdd FILL
XFILL_3_NOR2X1_126 gnd vdd FILL
XFILL_17_DFFSR_141 gnd vdd FILL
XFILL_58_DFFSR_97 gnd vdd FILL
XFILL_17_DFFSR_152 gnd vdd FILL
XFILL_3_NOR2X1_137 gnd vdd FILL
XFILL_17_DFFSR_1 gnd vdd FILL
XFILL_3_NOR2X1_148 gnd vdd FILL
XFILL_3_NOR2X1_159 gnd vdd FILL
XFILL_17_DFFSR_163 gnd vdd FILL
XFILL_17_DFFSR_174 gnd vdd FILL
XFILL_3_NOR2X1_7 gnd vdd FILL
XFILL_74_DFFSR_2 gnd vdd FILL
XFILL_6_CLKBUF1_6 gnd vdd FILL
XFILL_17_DFFSR_185 gnd vdd FILL
XFILL_17_DFFSR_196 gnd vdd FILL
XFILL_27_DFFSR_30 gnd vdd FILL
XFILL_27_DFFSR_41 gnd vdd FILL
XFILL_27_DFFSR_52 gnd vdd FILL
XFILL_27_DFFSR_63 gnd vdd FILL
XFILL_2_BUFX4_101 gnd vdd FILL
XFILL_27_DFFSR_74 gnd vdd FILL
XFILL_55_7_0 gnd vdd FILL
XFILL_27_DFFSR_85 gnd vdd FILL
XFILL_27_DFFSR_96 gnd vdd FILL
XFILL_27_4_2 gnd vdd FILL
XFILL_2_4_2 gnd vdd FILL
XFILL_13_NOR3X1_20 gnd vdd FILL
XFILL_13_NOR3X1_31 gnd vdd FILL
XFILL_67_DFFSR_40 gnd vdd FILL
XFILL_2_MUX2X1_5 gnd vdd FILL
XFILL_13_NOR3X1_42 gnd vdd FILL
XFILL_67_DFFSR_51 gnd vdd FILL
XFILL_20_MUX2X1_106 gnd vdd FILL
XFILL_20_MUX2X1_117 gnd vdd FILL
XFILL_63_DFFSR_220 gnd vdd FILL
XFILL_67_DFFSR_62 gnd vdd FILL
XFILL_20_MUX2X1_128 gnd vdd FILL
XFILL_6_BUFX4_100 gnd vdd FILL
XFILL_67_DFFSR_73 gnd vdd FILL
XFILL_20_MUX2X1_139 gnd vdd FILL
XFILL_63_DFFSR_231 gnd vdd FILL
XFILL_67_DFFSR_84 gnd vdd FILL
XFILL_63_DFFSR_242 gnd vdd FILL
XFILL_67_DFFSR_95 gnd vdd FILL
XFILL_63_DFFSR_253 gnd vdd FILL
XFILL_63_DFFSR_264 gnd vdd FILL
XFILL_63_DFFSR_275 gnd vdd FILL
XFILL_17_NOR3X1_30 gnd vdd FILL
XFILL_17_NOR3X1_41 gnd vdd FILL
XFILL_39_DFFSR_5 gnd vdd FILL
XFILL_17_NOR3X1_52 gnd vdd FILL
XFILL_8_NOR2X1_204 gnd vdd FILL
XFILL_67_DFFSR_230 gnd vdd FILL
XFILL_0_OAI22X1_13 gnd vdd FILL
XFILL_67_DFFSR_241 gnd vdd FILL
XFILL_0_OAI22X1_24 gnd vdd FILL
XFILL_0_OAI22X1_35 gnd vdd FILL
XFILL_67_DFFSR_252 gnd vdd FILL
XFILL_36_DFFSR_50 gnd vdd FILL
XFILL_0_OAI22X1_46 gnd vdd FILL
XFILL_10_3_2 gnd vdd FILL
XFILL_36_DFFSR_61 gnd vdd FILL
XFILL_67_DFFSR_263 gnd vdd FILL
XFILL_67_DFFSR_274 gnd vdd FILL
XFILL_22_CLKBUF1_4 gnd vdd FILL
XFILL_4_OAI21X1_15 gnd vdd FILL
XFILL_36_DFFSR_72 gnd vdd FILL
XFILL_36_DFFSR_83 gnd vdd FILL
XFILL_4_OAI21X1_26 gnd vdd FILL
XFILL_4_OAI21X1_37 gnd vdd FILL
XFILL_36_DFFSR_94 gnd vdd FILL
XFILL_0_NOR2X1_14 gnd vdd FILL
XFILL_0_NOR2X1_25 gnd vdd FILL
XFILL_4_OAI21X1_48 gnd vdd FILL
XAOI21X1_40 BUFX4_65/Y NOR2X1_202/B NOR2X1_200/Y gnd DFFSR_7/D vdd AOI21X1
XFILL_0_NOR2X1_36 gnd vdd FILL
XAOI21X1_51 BUFX4_97/Y NOR2X1_9/B NOR2X1_9/Y gnd DFFSR_270/D vdd AOI21X1
XFILL_0_NOR2X1_47 gnd vdd FILL
XAOI21X1_62 OAI21X1_45/Y NAND3X1_39/B DFFSR_1/D gnd AND2X2_3/B vdd AOI21X1
XFILL_0_NOR2X1_58 gnd vdd FILL
XAOI21X1_73 DFFSR_9/Q NOR2X1_52/Y NOR2X1_102/Y gnd NAND3X1_17/C vdd AOI21X1
XFILL_0_NOR2X1_69 gnd vdd FILL
XFILL_76_DFFSR_60 gnd vdd FILL
XFILL_26_CLKBUF1_3 gnd vdd FILL
XFILL_76_DFFSR_71 gnd vdd FILL
XFILL_76_DFFSR_82 gnd vdd FILL
XFILL_4_NOR2X1_13 gnd vdd FILL
XOAI21X1_2 OAI21X1_2/A OAI21X1_2/B OAI21X1_2/C gnd OAI21X1_2/Y vdd OAI21X1
XFILL_76_DFFSR_93 gnd vdd FILL
XFILL_45_DFFSR_209 gnd vdd FILL
XFILL_11_BUFX4_1 gnd vdd FILL
XFILL_4_NOR2X1_24 gnd vdd FILL
XFILL_3_NAND2X1_80 gnd vdd FILL
XFILL_4_NOR2X1_35 gnd vdd FILL
XFILL_4_NOR2X1_46 gnd vdd FILL
XFILL_3_NAND2X1_91 gnd vdd FILL
XFILL_4_NOR2X1_57 gnd vdd FILL
XFILL_9_0_1 gnd vdd FILL
XFILL_4_NOR2X1_68 gnd vdd FILL
XFILL_4_NOR2X1_79 gnd vdd FILL
XFILL_11_CLKBUF1_11 gnd vdd FILL
XFILL_16_NOR3X1_1 gnd vdd FILL
XFILL_8_NOR2X1_12 gnd vdd FILL
XFILL_11_CLKBUF1_22 gnd vdd FILL
XFILL_72_DFFSR_109 gnd vdd FILL
XFILL_49_DFFSR_208 gnd vdd FILL
XFILL_49_DFFSR_219 gnd vdd FILL
XFILL_11_CLKBUF1_33 gnd vdd FILL
XFILL_8_NOR2X1_23 gnd vdd FILL
XFILL_45_DFFSR_70 gnd vdd FILL
XFILL_8_NOR2X1_34 gnd vdd FILL
XFILL_45_DFFSR_81 gnd vdd FILL
XFILL_8_NOR2X1_45 gnd vdd FILL
XFILL_8_NOR2X1_56 gnd vdd FILL
XFILL_12_OAI22X1_7 gnd vdd FILL
XFILL_45_DFFSR_92 gnd vdd FILL
XFILL_8_NOR2X1_67 gnd vdd FILL
XFILL_8_NOR2X1_78 gnd vdd FILL
XFILL_8_NOR2X1_89 gnd vdd FILL
XFILL_76_DFFSR_108 gnd vdd FILL
XFILL_46_7_0 gnd vdd FILL
XFILL_76_DFFSR_119 gnd vdd FILL
XFILL_18_4_2 gnd vdd FILL
XFILL_85_DFFSR_80 gnd vdd FILL
XFILL_16_OAI22X1_6 gnd vdd FILL
XFILL_85_DFFSR_91 gnd vdd FILL
XFILL_14_DFFSR_80 gnd vdd FILL
XFILL_14_DFFSR_91 gnd vdd FILL
XFILL_60_2_2 gnd vdd FILL
XFILL_26_7 gnd vdd FILL
XFILL_30_DFFSR_220 gnd vdd FILL
XFILL_30_DFFSR_231 gnd vdd FILL
XFILL_30_DFFSR_242 gnd vdd FILL
XFILL_30_DFFSR_253 gnd vdd FILL
XFILL_30_DFFSR_264 gnd vdd FILL
XFILL_30_DFFSR_275 gnd vdd FILL
XFILL_54_DFFSR_90 gnd vdd FILL
XFILL_7_AOI21X1_80 gnd vdd FILL
XFILL_34_DFFSR_230 gnd vdd FILL
XFILL_34_DFFSR_241 gnd vdd FILL
XFILL_11_INVX4_1 gnd vdd FILL
XFILL_34_DFFSR_252 gnd vdd FILL
XFILL_34_DFFSR_263 gnd vdd FILL
XFILL_34_DFFSR_274 gnd vdd FILL
XFILL_0_MUX2X1_10 gnd vdd FILL
XFILL_0_MUX2X1_21 gnd vdd FILL
XFILL_1_INVX8_1 gnd vdd FILL
XFILL_0_MUX2X1_32 gnd vdd FILL
XFILL_0_MUX2X1_43 gnd vdd FILL
XFILL_0_MUX2X1_54 gnd vdd FILL
XFILL_61_DFFSR_130 gnd vdd FILL
XFILL_0_MUX2X1_65 gnd vdd FILL
XFILL_61_DFFSR_141 gnd vdd FILL
XFILL_61_DFFSR_152 gnd vdd FILL
XFILL_0_MUX2X1_76 gnd vdd FILL
XFILL_38_DFFSR_240 gnd vdd FILL
XFILL_0_MUX2X1_87 gnd vdd FILL
XFILL_38_DFFSR_251 gnd vdd FILL
XFILL_38_DFFSR_262 gnd vdd FILL
XFILL_61_DFFSR_163 gnd vdd FILL
XFILL_0_MUX2X1_98 gnd vdd FILL
XFILL_61_DFFSR_174 gnd vdd FILL
XFILL_38_DFFSR_273 gnd vdd FILL
XFILL_4_MUX2X1_20 gnd vdd FILL
XFILL_61_DFFSR_185 gnd vdd FILL
XFILL_4_MUX2X1_31 gnd vdd FILL
XFILL_61_DFFSR_196 gnd vdd FILL
XFILL_4_MUX2X1_42 gnd vdd FILL
XFILL_12_DFFSR_209 gnd vdd FILL
XFILL_4_MUX2X1_53 gnd vdd FILL
XFILL_4_MUX2X1_64 gnd vdd FILL
XFILL_65_DFFSR_140 gnd vdd FILL
XFILL_4_MUX2X1_75 gnd vdd FILL
XFILL_65_DFFSR_151 gnd vdd FILL
XFILL_10_OAI21X1_40 gnd vdd FILL
XFILL_65_DFFSR_162 gnd vdd FILL
XFILL_4_MUX2X1_86 gnd vdd FILL
XFILL_4_MUX2X1_97 gnd vdd FILL
XFILL_65_DFFSR_173 gnd vdd FILL
XFILL_65_DFFSR_184 gnd vdd FILL
XFILL_8_MUX2X1_30 gnd vdd FILL
XFILL_65_DFFSR_195 gnd vdd FILL
XFILL_16_DFFSR_208 gnd vdd FILL
XFILL_10_BUFX4_18 gnd vdd FILL
XFILL_8_MUX2X1_41 gnd vdd FILL
XFILL_16_DFFSR_219 gnd vdd FILL
XFILL_8_MUX2X1_52 gnd vdd FILL
XFILL_10_BUFX4_29 gnd vdd FILL
XFILL_13_NAND3X1_8 gnd vdd FILL
XFILL_8_MUX2X1_63 gnd vdd FILL
XFILL_69_DFFSR_150 gnd vdd FILL
XFILL_8_MUX2X1_74 gnd vdd FILL
XFILL_69_DFFSR_161 gnd vdd FILL
XFILL_6_DFFSR_90 gnd vdd FILL
XFILL_8_MUX2X1_85 gnd vdd FILL
XFILL_8_MUX2X1_96 gnd vdd FILL
XFILL_69_DFFSR_172 gnd vdd FILL
XFILL_37_7_0 gnd vdd FILL
XFILL_69_DFFSR_183 gnd vdd FILL
XFILL_69_DFFSR_194 gnd vdd FILL
XFILL_43_DFFSR_108 gnd vdd FILL
XFILL_43_DFFSR_119 gnd vdd FILL
XFILL_51_2_2 gnd vdd FILL
XFILL_47_DFFSR_107 gnd vdd FILL
XFILL_40_DFFSR_5 gnd vdd FILL
XFILL_47_DFFSR_118 gnd vdd FILL
XFILL_8_DFFSR_4 gnd vdd FILL
XFILL_20_MUX2X1_40 gnd vdd FILL
XFILL_47_DFFSR_129 gnd vdd FILL
XFILL_20_MUX2X1_51 gnd vdd FILL
XFILL_12_NAND3X1_16 gnd vdd FILL
XFILL_20_MUX2X1_62 gnd vdd FILL
XFILL_12_NAND3X1_27 gnd vdd FILL
XFILL_78_DFFSR_3 gnd vdd FILL
XFILL_20_MUX2X1_73 gnd vdd FILL
XFILL_20_6_0 gnd vdd FILL
XFILL_20_MUX2X1_84 gnd vdd FILL
XFILL_12_NAND3X1_38 gnd vdd FILL
XFILL_4_INVX1_19 gnd vdd FILL
XFILL_20_MUX2X1_95 gnd vdd FILL
XFILL_12_NAND3X1_49 gnd vdd FILL
XFILL_32_CLKBUF1_16 gnd vdd FILL
XFILL_32_CLKBUF1_27 gnd vdd FILL
XFILL_32_CLKBUF1_38 gnd vdd FILL
XFILL_2_BUFX4_17 gnd vdd FILL
XFILL_62_DFFSR_9 gnd vdd FILL
XFILL_2_BUFX4_28 gnd vdd FILL
XFILL_2_BUFX4_39 gnd vdd FILL
XFILL_59_3_2 gnd vdd FILL
XFILL_32_DFFSR_140 gnd vdd FILL
XFILL_32_DFFSR_151 gnd vdd FILL
XFILL_32_DFFSR_162 gnd vdd FILL
XFILL_32_DFFSR_173 gnd vdd FILL
XFILL_32_DFFSR_184 gnd vdd FILL
XFILL_32_DFFSR_195 gnd vdd FILL
XFILL_2_NAND3X1_11 gnd vdd FILL
XFILL_28_7_0 gnd vdd FILL
XFILL_2_NAND3X1_22 gnd vdd FILL
XFILL_3_7_0 gnd vdd FILL
XFILL_2_NAND3X1_33 gnd vdd FILL
XFILL_36_DFFSR_150 gnd vdd FILL
XFILL_2_NAND3X1_44 gnd vdd FILL
XFILL_36_DFFSR_161 gnd vdd FILL
XFILL_2_NAND3X1_55 gnd vdd FILL
XFILL_6_NAND2X1_13 gnd vdd FILL
XFILL_2_NAND3X1_66 gnd vdd FILL
XFILL_36_DFFSR_172 gnd vdd FILL
XFILL_6_NAND2X1_24 gnd vdd FILL
XFILL_2_NAND3X1_77 gnd vdd FILL
XFILL_36_DFFSR_183 gnd vdd FILL
XFILL_2_BUFX4_4 gnd vdd FILL
XFILL_2_NAND3X1_88 gnd vdd FILL
XFILL_36_DFFSR_194 gnd vdd FILL
XFILL_6_NAND2X1_35 gnd vdd FILL
XFILL_10_DFFSR_108 gnd vdd FILL
XFILL_2_NAND3X1_99 gnd vdd FILL
XFILL_6_NAND2X1_46 gnd vdd FILL
XFILL_6_NAND2X1_57 gnd vdd FILL
XFILL_10_DFFSR_119 gnd vdd FILL
XFILL_15_BUFX4_2 gnd vdd FILL
XFILL_6_NAND2X1_68 gnd vdd FILL
XFILL_6_NAND2X1_79 gnd vdd FILL
XFILL_42_2_2 gnd vdd FILL
XFILL_28_DFFSR_19 gnd vdd FILL
XMUX2X1_6 MUX2X1_6/A MUX2X1_6/B MUX2X1_7/S gnd MUX2X1_6/Y vdd MUX2X1
XFILL_14_DFFSR_107 gnd vdd FILL
XFILL_14_DFFSR_118 gnd vdd FILL
XFILL_11_6_0 gnd vdd FILL
XFILL_14_DFFSR_129 gnd vdd FILL
XFILL_68_DFFSR_18 gnd vdd FILL
XFILL_68_DFFSR_29 gnd vdd FILL
XFILL_82_DFFSR_240 gnd vdd FILL
XFILL_82_DFFSR_251 gnd vdd FILL
XFILL_82_DFFSR_262 gnd vdd FILL
XFILL_18_DFFSR_106 gnd vdd FILL
XFILL_82_DFFSR_273 gnd vdd FILL
XFILL_18_DFFSR_117 gnd vdd FILL
XFILL_18_DFFSR_128 gnd vdd FILL
XFILL_1_INVX1_8 gnd vdd FILL
XFILL_18_DFFSR_139 gnd vdd FILL
XFILL_13_AOI21X1_2 gnd vdd FILL
XCLKBUF1_7 BUFX4_9/Y gnd CLKBUF1_7/Y vdd CLKBUF1
XFILL_86_DFFSR_250 gnd vdd FILL
XFILL_6_AOI22X1_11 gnd vdd FILL
XFILL_10_NOR3X1_19 gnd vdd FILL
XFILL_86_DFFSR_261 gnd vdd FILL
XFILL_86_DFFSR_272 gnd vdd FILL
XFILL_37_DFFSR_17 gnd vdd FILL
XFILL_37_DFFSR_28 gnd vdd FILL
XFILL_37_DFFSR_39 gnd vdd FILL
XFILL_60_DFFSR_208 gnd vdd FILL
XFILL_60_DFFSR_219 gnd vdd FILL
XFILL_14_NOR3X1_18 gnd vdd FILL
XFILL_77_DFFSR_16 gnd vdd FILL
XFILL_14_NOR3X1_29 gnd vdd FILL
XFILL_21_CLKBUF1_12 gnd vdd FILL
XFILL_77_DFFSR_27 gnd vdd FILL
XFILL_77_DFFSR_38 gnd vdd FILL
XFILL_64_DFFSR_207 gnd vdd FILL
XFILL_21_CLKBUF1_23 gnd vdd FILL
XFILL_77_DFFSR_49 gnd vdd FILL
XBUFX4_101 INVX8_3/Y gnd MUX2X1_66/A vdd BUFX4
XFILL_21_CLKBUF1_34 gnd vdd FILL
XFILL_64_DFFSR_218 gnd vdd FILL
XFILL_64_DFFSR_229 gnd vdd FILL
XFILL_0_INVX1_12 gnd vdd FILL
XFILL_0_INVX1_23 gnd vdd FILL
XFILL_19_7_0 gnd vdd FILL
XFILL_0_INVX1_34 gnd vdd FILL
XFILL_4_CLKBUF1_16 gnd vdd FILL
XFILL_18_NOR3X1_17 gnd vdd FILL
XFILL_18_NOR3X1_28 gnd vdd FILL
XFILL_0_INVX1_45 gnd vdd FILL
XFILL_4_CLKBUF1_27 gnd vdd FILL
XFILL_1_AND2X2_4 gnd vdd FILL
XFILL_5_INVX8_2 gnd vdd FILL
XFILL_18_NOR3X1_39 gnd vdd FILL
XFILL_4_CLKBUF1_38 gnd vdd FILL
XNOR2X1_205 DFFSR_5/Q MUX2X1_22/S gnd NOR2X1_205/Y vdd NOR2X1
XFILL_0_INVX1_56 gnd vdd FILL
XFILL_68_DFFSR_206 gnd vdd FILL
XFILL_0_INVX1_67 gnd vdd FILL
XFILL_68_DFFSR_217 gnd vdd FILL
XFILL_0_INVX1_78 gnd vdd FILL
XFILL_46_DFFSR_15 gnd vdd FILL
XFILL_0_INVX1_89 gnd vdd FILL
XFILL_68_DFFSR_228 gnd vdd FILL
XFILL_46_DFFSR_26 gnd vdd FILL
XFILL_46_DFFSR_37 gnd vdd FILL
XFILL_68_DFFSR_239 gnd vdd FILL
XFILL_31_5 gnd vdd FILL
XFILL_46_DFFSR_48 gnd vdd FILL
XFILL_61_5_0 gnd vdd FILL
XFILL_46_DFFSR_59 gnd vdd FILL
XFILL_33_2_2 gnd vdd FILL
XFILL_2_NOR2X1_101 gnd vdd FILL
XFILL_24_4 gnd vdd FILL
XFILL_2_NOR2X1_112 gnd vdd FILL
XFILL_13_OAI21X1_17 gnd vdd FILL
XFILL_86_DFFSR_14 gnd vdd FILL
XFILL_13_OAI21X1_28 gnd vdd FILL
XFILL_2_NOR2X1_123 gnd vdd FILL
XFILL_86_DFFSR_25 gnd vdd FILL
XFILL_2_NOR2X1_134 gnd vdd FILL
XFILL_13_OAI21X1_39 gnd vdd FILL
XFILL_22_DFFSR_2 gnd vdd FILL
XFILL_2_NOR2X1_145 gnd vdd FILL
XFILL_86_DFFSR_36 gnd vdd FILL
XFILL_17_3 gnd vdd FILL
XFILL_2_NOR2X1_156 gnd vdd FILL
XFILL_86_DFFSR_47 gnd vdd FILL
XFILL_86_DFFSR_58 gnd vdd FILL
XFILL_15_DFFSR_14 gnd vdd FILL
XFILL_2_NOR2X1_167 gnd vdd FILL
XFILL_86_DFFSR_69 gnd vdd FILL
XFILL_15_DFFSR_25 gnd vdd FILL
XFILL_2_NOR2X1_178 gnd vdd FILL
XFILL_15_DFFSR_36 gnd vdd FILL
XFILL_2_NOR2X1_189 gnd vdd FILL
XFILL_15_DFFSR_47 gnd vdd FILL
XFILL_15_DFFSR_58 gnd vdd FILL
XFILL_26_14 gnd vdd FILL
XFILL_15_DFFSR_69 gnd vdd FILL
XFILL_55_DFFSR_13 gnd vdd FILL
XFILL_55_DFFSR_24 gnd vdd FILL
XFILL_55_DFFSR_35 gnd vdd FILL
XFILL_55_DFFSR_46 gnd vdd FILL
XFILL_55_DFFSR_57 gnd vdd FILL
XFILL_55_DFFSR_68 gnd vdd FILL
XFILL_55_DFFSR_79 gnd vdd FILL
XFILL_53_DFFSR_250 gnd vdd FILL
XFILL_53_DFFSR_261 gnd vdd FILL
XFILL_53_DFFSR_272 gnd vdd FILL
XFILL_2_MUX2X1_107 gnd vdd FILL
XFILL_2_MUX2X1_118 gnd vdd FILL
XFILL_2_MUX2X1_129 gnd vdd FILL
XFILL_44_DFFSR_6 gnd vdd FILL
XFILL_24_DFFSR_12 gnd vdd FILL
XFILL_7_NOR2X1_201 gnd vdd FILL
XFILL_24_DFFSR_23 gnd vdd FILL
XFILL_24_DFFSR_34 gnd vdd FILL
XFILL_24_DFFSR_45 gnd vdd FILL
XFILL_80_DFFSR_150 gnd vdd FILL
XFILL_24_DFFSR_56 gnd vdd FILL
XFILL_80_DFFSR_161 gnd vdd FILL
XFILL_24_DFFSR_67 gnd vdd FILL
XFILL_57_DFFSR_260 gnd vdd FILL
XFILL_57_DFFSR_271 gnd vdd FILL
XFILL_24_DFFSR_78 gnd vdd FILL
XFILL_12_CLKBUF1_1 gnd vdd FILL
XFILL_80_DFFSR_172 gnd vdd FILL
XFILL_24_DFFSR_89 gnd vdd FILL
XFILL_80_DFFSR_183 gnd vdd FILL
XFILL_3_OAI21X1_12 gnd vdd FILL
XFILL_80_DFFSR_194 gnd vdd FILL
XFILL_3_OAI21X1_23 gnd vdd FILL
XFILL_31_DFFSR_207 gnd vdd FILL
XFILL_64_DFFSR_11 gnd vdd FILL
XFILL_0_DFFSR_220 gnd vdd FILL
XFILL_3_OAI21X1_34 gnd vdd FILL
XFILL_64_DFFSR_22 gnd vdd FILL
XFILL_31_DFFSR_218 gnd vdd FILL
XFILL_3_OAI21X1_45 gnd vdd FILL
XFILL_64_DFFSR_33 gnd vdd FILL
XFILL_0_DFFSR_231 gnd vdd FILL
XFILL_0_DFFSR_242 gnd vdd FILL
XFILL_31_DFFSR_229 gnd vdd FILL
XFILL_64_DFFSR_44 gnd vdd FILL
XFILL_64_DFFSR_55 gnd vdd FILL
XFILL_0_DFFSR_253 gnd vdd FILL
XFILL_84_DFFSR_160 gnd vdd FILL
XFILL_0_DFFSR_264 gnd vdd FILL
XFILL_0_DFFSR_275 gnd vdd FILL
XFILL_64_DFFSR_66 gnd vdd FILL
XFILL_64_DFFSR_77 gnd vdd FILL
XFILL_84_DFFSR_171 gnd vdd FILL
XFILL_64_DFFSR_88 gnd vdd FILL
XFILL_84_DFFSR_182 gnd vdd FILL
XFILL_64_DFFSR_99 gnd vdd FILL
XFILL_84_DFFSR_193 gnd vdd FILL
XFILL_35_DFFSR_206 gnd vdd FILL
XFILL_52_5_0 gnd vdd FILL
XFILL_35_DFFSR_217 gnd vdd FILL
XFILL_4_DFFSR_230 gnd vdd FILL
XFILL_7_DFFSR_13 gnd vdd FILL
XFILL_35_DFFSR_228 gnd vdd FILL
XFILL_24_2_2 gnd vdd FILL
XFILL_7_DFFSR_24 gnd vdd FILL
XFILL_4_DFFSR_241 gnd vdd FILL
XFILL_7_DFFSR_35 gnd vdd FILL
XFILL_35_DFFSR_239 gnd vdd FILL
XFILL_4_DFFSR_252 gnd vdd FILL
XFILL_33_DFFSR_10 gnd vdd FILL
XFILL_7_DFFSR_46 gnd vdd FILL
XFILL_4_DFFSR_263 gnd vdd FILL
XFILL_4_DFFSR_274 gnd vdd FILL
XFILL_33_DFFSR_21 gnd vdd FILL
XFILL_7_DFFSR_57 gnd vdd FILL
XFILL_33_DFFSR_32 gnd vdd FILL
XFILL_33_DFFSR_43 gnd vdd FILL
XFILL_7_DFFSR_68 gnd vdd FILL
XFILL_1_MUX2X1_19 gnd vdd FILL
XFILL_62_DFFSR_106 gnd vdd FILL
XFILL_7_DFFSR_79 gnd vdd FILL
XFILL_33_DFFSR_54 gnd vdd FILL
XFILL_39_DFFSR_205 gnd vdd FILL
XFILL_33_DFFSR_65 gnd vdd FILL
XFILL_10_CLKBUF1_30 gnd vdd FILL
XFILL_39_DFFSR_216 gnd vdd FILL
XFILL_62_DFFSR_117 gnd vdd FILL
XFILL_10_CLKBUF1_41 gnd vdd FILL
XFILL_33_DFFSR_76 gnd vdd FILL
XFILL_39_DFFSR_227 gnd vdd FILL
XFILL_8_DFFSR_240 gnd vdd FILL
XFILL_62_DFFSR_128 gnd vdd FILL
XFILL_33_DFFSR_87 gnd vdd FILL
XFILL_62_DFFSR_139 gnd vdd FILL
XFILL_33_DFFSR_98 gnd vdd FILL
XFILL_8_DFFSR_251 gnd vdd FILL
XFILL_39_DFFSR_238 gnd vdd FILL
XFILL_39_DFFSR_249 gnd vdd FILL
XFILL_8_DFFSR_262 gnd vdd FILL
XFILL_73_DFFSR_20 gnd vdd FILL
XFILL_8_DFFSR_273 gnd vdd FILL
XFILL_73_DFFSR_31 gnd vdd FILL
XFILL_5_MUX2X1_18 gnd vdd FILL
XFILL_73_DFFSR_42 gnd vdd FILL
XFILL_66_DFFSR_105 gnd vdd FILL
XFILL_5_MUX2X1_29 gnd vdd FILL
XFILL_73_DFFSR_53 gnd vdd FILL
XFILL_73_DFFSR_64 gnd vdd FILL
XFILL_66_DFFSR_116 gnd vdd FILL
XFILL_73_DFFSR_75 gnd vdd FILL
XFILL_66_DFFSR_127 gnd vdd FILL
XFILL_66_DFFSR_138 gnd vdd FILL
XFILL_73_DFFSR_86 gnd vdd FILL
XFILL_66_DFFSR_149 gnd vdd FILL
XFILL_73_DFFSR_97 gnd vdd FILL
XFILL_9_MUX2X1_17 gnd vdd FILL
XFILL_9_MUX2X1_28 gnd vdd FILL
XFILL_6_BUFX4_5 gnd vdd FILL
XFILL_9_MUX2X1_39 gnd vdd FILL
XFILL_42_DFFSR_30 gnd vdd FILL
XFILL_19_MUX2X1_110 gnd vdd FILL
XFILL_13_NOR3X1_5 gnd vdd FILL
XFILL_1_AOI22X1_2 gnd vdd FILL
XFILL_42_DFFSR_41 gnd vdd FILL
XFILL_19_MUX2X1_121 gnd vdd FILL
XFILL_13_OAI21X1_5 gnd vdd FILL
XFILL_10_NOR2X1_30 gnd vdd FILL
XFILL_42_DFFSR_52 gnd vdd FILL
XFILL_42_DFFSR_63 gnd vdd FILL
XFILL_10_NOR2X1_41 gnd vdd FILL
XFILL_19_MUX2X1_132 gnd vdd FILL
XFILL_10_NOR2X1_52 gnd vdd FILL
XFILL_42_DFFSR_74 gnd vdd FILL
XFILL_19_MUX2X1_143 gnd vdd FILL
XFILL_20_DFFSR_250 gnd vdd FILL
XFILL_19_MUX2X1_154 gnd vdd FILL
XFILL_42_DFFSR_85 gnd vdd FILL
XFILL_10_NOR2X1_63 gnd vdd FILL
XFILL_20_DFFSR_261 gnd vdd FILL
XFILL_19_MUX2X1_165 gnd vdd FILL
XFILL_20_DFFSR_272 gnd vdd FILL
XFILL_10_NOR2X1_74 gnd vdd FILL
XFILL_7_3_2 gnd vdd FILL
XFILL_42_DFFSR_96 gnd vdd FILL
XFILL_1_INVX1_201 gnd vdd FILL
XBUFX4_18 rst_n gnd BUFX4_47/A vdd BUFX4
XFILL_1_INVX1_212 gnd vdd FILL
XFILL_10_NOR2X1_85 gnd vdd FILL
XFILL_19_MUX2X1_176 gnd vdd FILL
XFILL_19_MUX2X1_187 gnd vdd FILL
XBUFX4_29 rst_n gnd BUFX4_44/A vdd BUFX4
XFILL_1_INVX1_223 gnd vdd FILL
XFILL_10_NOR2X1_96 gnd vdd FILL
XFILL_82_DFFSR_40 gnd vdd FILL
XFILL_5_AOI22X1_1 gnd vdd FILL
XFILL_82_DFFSR_51 gnd vdd FILL
XFILL_82_DFFSR_62 gnd vdd FILL
XFILL_82_DFFSR_73 gnd vdd FILL
XFILL_82_DFFSR_84 gnd vdd FILL
XFILL_11_DFFSR_40 gnd vdd FILL
XFILL_24_DFFSR_260 gnd vdd FILL
XFILL_82_DFFSR_95 gnd vdd FILL
XFILL_24_DFFSR_271 gnd vdd FILL
XFILL_11_DFFSR_51 gnd vdd FILL
XFILL_5_INVX1_200 gnd vdd FILL
XFILL_21_MUX2X1_16 gnd vdd FILL
XFILL_11_DFFSR_62 gnd vdd FILL
XFILL_5_INVX1_211 gnd vdd FILL
XFILL_5_INVX1_9 gnd vdd FILL
XFILL_11_DFFSR_73 gnd vdd FILL
XFILL_21_MUX2X1_27 gnd vdd FILL
XFILL_5_INVX1_222 gnd vdd FILL
XFILL_11_DFFSR_84 gnd vdd FILL
XFILL_21_MUX2X1_38 gnd vdd FILL
XFILL_11_DFFSR_95 gnd vdd FILL
XFILL_21_MUX2X1_49 gnd vdd FILL
XFILL_51_DFFSR_160 gnd vdd FILL
XFILL_2_BUFX2_1 gnd vdd FILL
XFILL_22_NOR3X1_3 gnd vdd FILL
XFILL_43_5_0 gnd vdd FILL
XFILL_28_DFFSR_270 gnd vdd FILL
XFILL_51_DFFSR_171 gnd vdd FILL
XFILL_51_DFFSR_50 gnd vdd FILL
XFILL_15_2_2 gnd vdd FILL
XFILL_51_DFFSR_182 gnd vdd FILL
XFILL_51_DFFSR_193 gnd vdd FILL
XFILL_51_DFFSR_61 gnd vdd FILL
XFILL_51_DFFSR_72 gnd vdd FILL
XFILL_51_DFFSR_83 gnd vdd FILL
XFILL_51_DFFSR_94 gnd vdd FILL
XFILL_55_DFFSR_170 gnd vdd FILL
XFILL_55_DFFSR_181 gnd vdd FILL
XFILL_55_DFFSR_192 gnd vdd FILL
XFILL_20_DFFSR_60 gnd vdd FILL
XFILL_9_MUX2X1_160 gnd vdd FILL
XFILL_20_DFFSR_71 gnd vdd FILL
XFILL_20_DFFSR_82 gnd vdd FILL
XFILL_9_MUX2X1_171 gnd vdd FILL
XFILL_20_DFFSR_93 gnd vdd FILL
XFILL_9_MUX2X1_182 gnd vdd FILL
XFILL_59_DFFSR_180 gnd vdd FILL
XFILL_5_NOR3X1_4 gnd vdd FILL
XFILL_9_MUX2X1_193 gnd vdd FILL
XFILL_33_DFFSR_105 gnd vdd FILL
XFILL_59_DFFSR_191 gnd vdd FILL
XFILL_9_INVX8_3 gnd vdd FILL
XFILL_31_NOR3X1_1 gnd vdd FILL
XFILL_33_DFFSR_116 gnd vdd FILL
XFILL_10_NAND2X1_7 gnd vdd FILL
XFILL_2_DFFSR_140 gnd vdd FILL
XFILL_33_DFFSR_127 gnd vdd FILL
XFILL_33_DFFSR_138 gnd vdd FILL
XFILL_2_DFFSR_151 gnd vdd FILL
XFILL_2_DFFSR_162 gnd vdd FILL
XFILL_33_DFFSR_149 gnd vdd FILL
XFILL_60_DFFSR_70 gnd vdd FILL
XFILL_2_DFFSR_173 gnd vdd FILL
XFILL_60_DFFSR_81 gnd vdd FILL
XFILL_2_DFFSR_184 gnd vdd FILL
XFILL_60_DFFSR_92 gnd vdd FILL
XFILL_2_DFFSR_195 gnd vdd FILL
XFILL_37_DFFSR_104 gnd vdd FILL
XFILL_37_DFFSR_115 gnd vdd FILL
XFILL_37_DFFSR_126 gnd vdd FILL
XFILL_26_DFFSR_3 gnd vdd FILL
XFILL_37_DFFSR_137 gnd vdd FILL
XFILL_6_DFFSR_150 gnd vdd FILL
XFILL_6_DFFSR_161 gnd vdd FILL
XFILL_37_DFFSR_148 gnd vdd FILL
XFILL_11_NAND3X1_13 gnd vdd FILL
XFILL_3_DFFSR_50 gnd vdd FILL
XFILL_6_DFFSR_172 gnd vdd FILL
XFILL_37_DFFSR_159 gnd vdd FILL
XFILL_3_DFFSR_61 gnd vdd FILL
XFILL_11_NAND3X1_24 gnd vdd FILL
XFILL_83_DFFSR_4 gnd vdd FILL
XFILL_10_MUX2X1_70 gnd vdd FILL
XFILL_11_NAND3X1_35 gnd vdd FILL
XFILL_10_MUX2X1_81 gnd vdd FILL
XFILL_6_DFFSR_183 gnd vdd FILL
XFILL_3_DFFSR_72 gnd vdd FILL
XFILL_3_DFFSR_83 gnd vdd FILL
XFILL_10_MUX2X1_92 gnd vdd FILL
XFILL_6_DFFSR_194 gnd vdd FILL
XFILL_11_NAND3X1_46 gnd vdd FILL
XFILL_11_NAND3X1_57 gnd vdd FILL
XFILL_3_DFFSR_94 gnd vdd FILL
XFILL_11_NAND3X1_68 gnd vdd FILL
XFILL_31_CLKBUF1_13 gnd vdd FILL
XFILL_2_INVX2_1 gnd vdd FILL
XFILL_11_NAND3X1_79 gnd vdd FILL
XFILL_31_CLKBUF1_24 gnd vdd FILL
XFILL_31_CLKBUF1_35 gnd vdd FILL
XFILL_65_1_2 gnd vdd FILL
XFILL_14_MUX2X1_80 gnd vdd FILL
XFILL_14_MUX2X1_91 gnd vdd FILL
XFILL_2_NOR3X1_40 gnd vdd FILL
XFILL_2_NOR3X1_51 gnd vdd FILL
XFILL_83_DFFSR_205 gnd vdd FILL
XFILL_83_DFFSR_216 gnd vdd FILL
XFILL_34_5_0 gnd vdd FILL
XFILL_83_DFFSR_227 gnd vdd FILL
XFILL_10_DFFSR_9 gnd vdd FILL
XFILL_83_DFFSR_238 gnd vdd FILL
XFILL_83_DFFSR_249 gnd vdd FILL
XFILL_18_MUX2X1_90 gnd vdd FILL
XFILL_22_1 gnd vdd FILL
XFILL_6_NOR3X1_50 gnd vdd FILL
XFILL_48_DFFSR_7 gnd vdd FILL
XFILL_87_DFFSR_204 gnd vdd FILL
XFILL_87_DFFSR_215 gnd vdd FILL
XFILL_87_DFFSR_226 gnd vdd FILL
XFILL_87_DFFSR_237 gnd vdd FILL
XFILL_87_DFFSR_248 gnd vdd FILL
XFILL_22_DFFSR_170 gnd vdd FILL
XFILL_87_DFFSR_259 gnd vdd FILL
XFILL_3_INVX1_110 gnd vdd FILL
XFILL_22_DFFSR_181 gnd vdd FILL
XFILL_22_DFFSR_192 gnd vdd FILL
XFILL_3_INVX1_121 gnd vdd FILL
XFILL_3_INVX1_132 gnd vdd FILL
XFILL_3_INVX1_143 gnd vdd FILL
XFILL_3_INVX1_154 gnd vdd FILL
XFILL_1_NAND3X1_30 gnd vdd FILL
XFILL_3_INVX1_165 gnd vdd FILL
XFILL_1_NAND3X1_41 gnd vdd FILL
XFILL_1_NAND3X1_52 gnd vdd FILL
XFILL_5_NAND2X1_10 gnd vdd FILL
XFILL_3_INVX1_176 gnd vdd FILL
XFILL_3_INVX1_187 gnd vdd FILL
XFILL_5_NAND2X1_21 gnd vdd FILL
XFILL_1_NAND3X1_63 gnd vdd FILL
XFILL_26_DFFSR_180 gnd vdd FILL
XFILL_1_NAND3X1_74 gnd vdd FILL
XFILL_3_INVX1_198 gnd vdd FILL
XFILL_5_NAND2X1_32 gnd vdd FILL
XFILL_1_NAND3X1_85 gnd vdd FILL
XFILL_7_INVX1_120 gnd vdd FILL
XFILL_26_DFFSR_191 gnd vdd FILL
XFILL_1_NAND3X1_96 gnd vdd FILL
XFILL_5_NAND2X1_43 gnd vdd FILL
XFILL_7_INVX1_131 gnd vdd FILL
XFILL_5_NAND2X1_54 gnd vdd FILL
XFILL_5_NAND2X1_65 gnd vdd FILL
XFILL_7_INVX1_142 gnd vdd FILL
XFILL_7_INVX1_153 gnd vdd FILL
XFILL_5_NAND2X1_76 gnd vdd FILL
XFILL_7_INVX1_164 gnd vdd FILL
XFILL_5_NAND2X1_87 gnd vdd FILL
XFILL_7_INVX1_175 gnd vdd FILL
XFILL_7_INVX1_186 gnd vdd FILL
XFILL_7_INVX1_197 gnd vdd FILL
XFILL_13_CLKBUF1_18 gnd vdd FILL
XFILL_13_CLKBUF1_29 gnd vdd FILL
XFILL_1_OAI22X1_5 gnd vdd FILL
XFILL_56_1_2 gnd vdd FILL
XFILL_72_DFFSR_270 gnd vdd FILL
XFILL_11_NOR2X1_103 gnd vdd FILL
XFILL_5_OAI22X1_4 gnd vdd FILL
XFILL_11_NOR2X1_114 gnd vdd FILL
XFILL_11_NOR2X1_125 gnd vdd FILL
XFILL_11_NOR2X1_136 gnd vdd FILL
XFILL_11_NOR2X1_147 gnd vdd FILL
XFILL_25_5_0 gnd vdd FILL
XFILL_0_5_0 gnd vdd FILL
XFILL_11_NOR2X1_158 gnd vdd FILL
XFILL_11_NOR2X1_169 gnd vdd FILL
XFILL_50_DFFSR_205 gnd vdd FILL
XFILL_9_AOI21X1_10 gnd vdd FILL
XFILL_50_DFFSR_216 gnd vdd FILL
XFILL_9_AOI21X1_21 gnd vdd FILL
XFILL_9_OAI22X1_3 gnd vdd FILL
XFILL_9_AOI21X1_32 gnd vdd FILL
XFILL_50_DFFSR_227 gnd vdd FILL
XFILL_50_DFFSR_238 gnd vdd FILL
XFILL_9_AOI21X1_43 gnd vdd FILL
XFILL_50_DFFSR_249 gnd vdd FILL
XFILL_9_AOI21X1_54 gnd vdd FILL
XFILL_19_OAI22X1_12 gnd vdd FILL
XFILL_9_AOI21X1_65 gnd vdd FILL
XFILL_19_OAI22X1_23 gnd vdd FILL
XFILL_9_AOI21X1_76 gnd vdd FILL
XFILL_20_CLKBUF1_20 gnd vdd FILL
XFILL_19_OAI22X1_34 gnd vdd FILL
XFILL_54_DFFSR_204 gnd vdd FILL
XFILL_19_OAI22X1_45 gnd vdd FILL
XFILL_54_DFFSR_215 gnd vdd FILL
XFILL_20_CLKBUF1_31 gnd vdd FILL
XFILL_20_CLKBUF1_42 gnd vdd FILL
XFILL_54_DFFSR_226 gnd vdd FILL
XFILL_54_DFFSR_237 gnd vdd FILL
XFILL_54_DFFSR_248 gnd vdd FILL
XFILL_3_CLKBUF1_13 gnd vdd FILL
XFILL_54_DFFSR_259 gnd vdd FILL
XFILL_3_CLKBUF1_24 gnd vdd FILL
XFILL_3_CLKBUF1_35 gnd vdd FILL
XFILL_81_DFFSR_104 gnd vdd FILL
XFILL_11_MUX2X1_109 gnd vdd FILL
XFILL_58_DFFSR_203 gnd vdd FILL
XFILL_81_DFFSR_115 gnd vdd FILL
XFILL_58_DFFSR_214 gnd vdd FILL
XFILL_81_DFFSR_126 gnd vdd FILL
XFILL_58_DFFSR_225 gnd vdd FILL
XFILL_81_DFFSR_137 gnd vdd FILL
XFILL_58_DFFSR_236 gnd vdd FILL
XFILL_81_DFFSR_148 gnd vdd FILL
XFILL_6_BUFX2_2 gnd vdd FILL
XFILL_58_DFFSR_247 gnd vdd FILL
XFILL_81_DFFSR_159 gnd vdd FILL
XFILL_58_DFFSR_258 gnd vdd FILL
XFILL_58_DFFSR_269 gnd vdd FILL
XFILL_1_DFFSR_207 gnd vdd FILL
XFILL_85_DFFSR_103 gnd vdd FILL
XFILL_85_DFFSR_114 gnd vdd FILL
XFILL_1_DFFSR_218 gnd vdd FILL
XFILL_12_OAI21X1_14 gnd vdd FILL
XFILL_1_NOR2X1_120 gnd vdd FILL
XFILL_12_OAI21X1_25 gnd vdd FILL
XFILL_1_DFFSR_229 gnd vdd FILL
XFILL_85_DFFSR_125 gnd vdd FILL
XFILL_85_DFFSR_136 gnd vdd FILL
XFILL_8_6_0 gnd vdd FILL
XFILL_12_OAI21X1_36 gnd vdd FILL
XFILL_1_NOR2X1_131 gnd vdd FILL
XFILL_85_DFFSR_147 gnd vdd FILL
XFILL_1_NOR2X1_142 gnd vdd FILL
XFILL_85_DFFSR_158 gnd vdd FILL
XFILL_1_NOR2X1_153 gnd vdd FILL
XFILL_12_OAI21X1_47 gnd vdd FILL
XFILL_85_DFFSR_169 gnd vdd FILL
XFILL_1_NOR2X1_164 gnd vdd FILL
XFILL_17_CLKBUF1_9 gnd vdd FILL
XFILL_1_NOR2X1_175 gnd vdd FILL
XFILL_65_DFFSR_1 gnd vdd FILL
XFILL_5_DFFSR_206 gnd vdd FILL
XFILL_8_BUFX4_10 gnd vdd FILL
XFILL_1_NOR2X1_186 gnd vdd FILL
XFILL_5_DFFSR_217 gnd vdd FILL
XFILL_1_NOR2X1_197 gnd vdd FILL
XFILL_2_NAND3X1_6 gnd vdd FILL
XFILL_8_BUFX4_21 gnd vdd FILL
XFILL_5_DFFSR_228 gnd vdd FILL
XFILL_8_BUFX4_32 gnd vdd FILL
XFILL_47_1_2 gnd vdd FILL
XFILL_8_BUFX4_43 gnd vdd FILL
XFILL_5_DFFSR_239 gnd vdd FILL
XFILL_8_BUFX4_54 gnd vdd FILL
XFILL_43_DFFSR_19 gnd vdd FILL
XFILL_13_BUFX4_104 gnd vdd FILL
XFILL_8_BUFX4_65 gnd vdd FILL
XFILL_8_BUFX4_76 gnd vdd FILL
XFILL_11_NAND2X1_90 gnd vdd FILL
XFILL_9_OAI22X1_40 gnd vdd FILL
XFILL_8_BUFX4_87 gnd vdd FILL
XFILL_9_DFFSR_205 gnd vdd FILL
XFILL_9_OAI22X1_51 gnd vdd FILL
XFILL_6_NAND3X1_5 gnd vdd FILL
XFILL_8_BUFX4_98 gnd vdd FILL
XFILL_9_DFFSR_216 gnd vdd FILL
XFILL_9_DFFSR_227 gnd vdd FILL
XFILL_9_DFFSR_238 gnd vdd FILL
XFILL_16_5_0 gnd vdd FILL
XFILL_9_DFFSR_249 gnd vdd FILL
XFILL_83_DFFSR_18 gnd vdd FILL
XFILL_83_DFFSR_29 gnd vdd FILL
XFILL_1_MUX2X1_104 gnd vdd FILL
XFILL_1_MUX2X1_115 gnd vdd FILL
XNAND3X1_120 DFFSR_26/Q BUFX4_6/Y NOR2X1_38/Y gnd NAND3X1_126/A vdd NAND3X1
XNAND3X1_131 DFFSR_83/Q BUFX4_1/Y NOR2X1_44/Y gnd OAI21X1_24/C vdd NAND3X1
XFILL_1_MUX2X1_126 gnd vdd FILL
XFILL_12_DFFSR_18 gnd vdd FILL
XFILL_12_DFFSR_29 gnd vdd FILL
XFILL_1_MUX2X1_137 gnd vdd FILL
XFILL_1_MUX2X1_148 gnd vdd FILL
XFILL_1_MUX2X1_159 gnd vdd FILL
XFILL_30_0_2 gnd vdd FILL
XFILL_87_DFFSR_5 gnd vdd FILL
XFILL_70_DFFSR_180 gnd vdd FILL
XFILL_6_INVX2_2 gnd vdd FILL
XFILL_2_OAI21X1_20 gnd vdd FILL
XFILL_52_DFFSR_17 gnd vdd FILL
XFILL_70_DFFSR_191 gnd vdd FILL
XFILL_2_OAI21X1_31 gnd vdd FILL
XFILL_52_DFFSR_28 gnd vdd FILL
XFILL_21_DFFSR_204 gnd vdd FILL
XFILL_21_DFFSR_215 gnd vdd FILL
XFILL_52_DFFSR_39 gnd vdd FILL
XFILL_2_OAI21X1_42 gnd vdd FILL
XFILL_21_DFFSR_226 gnd vdd FILL
XFILL_11_NOR2X1_17 gnd vdd FILL
XFILL_11_NOR2X1_28 gnd vdd FILL
XFILL_21_DFFSR_237 gnd vdd FILL
XFILL_11_NOR2X1_39 gnd vdd FILL
XFILL_21_DFFSR_248 gnd vdd FILL
XFILL_21_DFFSR_259 gnd vdd FILL
XFILL_74_DFFSR_190 gnd vdd FILL
XFILL_25_DFFSR_203 gnd vdd FILL
XFILL_9_MUX2X1_9 gnd vdd FILL
XFILL_25_DFFSR_214 gnd vdd FILL
XFILL_25_DFFSR_225 gnd vdd FILL
XFILL_21_DFFSR_16 gnd vdd FILL
XFILL_25_DFFSR_236 gnd vdd FILL
XFILL_25_DFFSR_247 gnd vdd FILL
XFILL_21_DFFSR_27 gnd vdd FILL
XFILL_21_DFFSR_38 gnd vdd FILL
XFILL_25_DFFSR_258 gnd vdd FILL
XFILL_25_DFFSR_269 gnd vdd FILL
XFILL_12_BUFX4_70 gnd vdd FILL
XFILL_21_DFFSR_49 gnd vdd FILL
XFILL_12_BUFX4_81 gnd vdd FILL
XFILL_6_INVX1_209 gnd vdd FILL
XFILL_52_DFFSR_103 gnd vdd FILL
XFILL_29_DFFSR_202 gnd vdd FILL
XFILL_12_BUFX4_92 gnd vdd FILL
XFILL_29_DFFSR_213 gnd vdd FILL
XFILL_52_DFFSR_114 gnd vdd FILL
XFILL_29_DFFSR_224 gnd vdd FILL
XFILL_52_DFFSR_125 gnd vdd FILL
XFILL_52_DFFSR_136 gnd vdd FILL
XFILL_29_DFFSR_235 gnd vdd FILL
XFILL_61_DFFSR_15 gnd vdd FILL
XFILL_52_DFFSR_147 gnd vdd FILL
XFILL_52_DFFSR_158 gnd vdd FILL
XFILL_61_DFFSR_26 gnd vdd FILL
XFILL_29_DFFSR_246 gnd vdd FILL
XFILL_61_DFFSR_37 gnd vdd FILL
XFILL_29_DFFSR_257 gnd vdd FILL
XFILL_66_4_0 gnd vdd FILL
XFILL_29_DFFSR_268 gnd vdd FILL
XFILL_52_DFFSR_169 gnd vdd FILL
XFILL_61_DFFSR_48 gnd vdd FILL
XFILL_61_DFFSR_59 gnd vdd FILL
XFILL_56_DFFSR_102 gnd vdd FILL
XFILL_38_1_2 gnd vdd FILL
XFILL_56_DFFSR_113 gnd vdd FILL
XFILL_56_DFFSR_124 gnd vdd FILL
XFILL_4_NAND3X1_18 gnd vdd FILL
XFILL_56_DFFSR_135 gnd vdd FILL
XFILL_4_NAND3X1_29 gnd vdd FILL
XFILL_56_DFFSR_146 gnd vdd FILL
XFILL_56_DFFSR_157 gnd vdd FILL
XFILL_4_DFFSR_17 gnd vdd FILL
XFILL_56_DFFSR_168 gnd vdd FILL
XFILL_4_DFFSR_28 gnd vdd FILL
XFILL_56_DFFSR_179 gnd vdd FILL
XFILL_30_DFFSR_14 gnd vdd FILL
XFILL_4_DFFSR_39 gnd vdd FILL
XFILL_30_DFFSR_25 gnd vdd FILL
XFILL_30_DFFSR_36 gnd vdd FILL
XFILL_30_DFFSR_47 gnd vdd FILL
XFILL_30_DFFSR_58 gnd vdd FILL
XFILL_6_INVX1_60 gnd vdd FILL
XFILL_30_DFFSR_69 gnd vdd FILL
XFILL_18_MUX2X1_140 gnd vdd FILL
XFILL_6_INVX1_71 gnd vdd FILL
XFILL_6_INVX1_82 gnd vdd FILL
XFILL_18_MUX2X1_151 gnd vdd FILL
XFILL_6_INVX1_93 gnd vdd FILL
XFILL_70_DFFSR_13 gnd vdd FILL
XFILL_18_MUX2X1_162 gnd vdd FILL
XFILL_3_DFFSR_105 gnd vdd FILL
XFILL_18_MUX2X1_173 gnd vdd FILL
XFILL_70_DFFSR_24 gnd vdd FILL
XFILL_21_0_2 gnd vdd FILL
XFILL_3_DFFSR_116 gnd vdd FILL
XFILL_70_DFFSR_35 gnd vdd FILL
XFILL_3_DFFSR_127 gnd vdd FILL
XFILL_18_MUX2X1_184 gnd vdd FILL
XFILL_3_DFFSR_138 gnd vdd FILL
XFILL_70_DFFSR_46 gnd vdd FILL
XFILL_13_MUX2X1_3 gnd vdd FILL
XFILL_3_DFFSR_149 gnd vdd FILL
XFILL_70_DFFSR_57 gnd vdd FILL
XFILL_70_DFFSR_68 gnd vdd FILL
XFILL_70_DFFSR_79 gnd vdd FILL
XFILL_7_DFFSR_104 gnd vdd FILL
XFILL_11_MUX2X1_13 gnd vdd FILL
XFILL_7_DFFSR_115 gnd vdd FILL
XDFFSR_140 DFFSR_140/Q CLKBUF1_8/Y DFFSR_58/R vdd DFFSR_140/D gnd vdd DFFSR
XFILL_7_DFFSR_126 gnd vdd FILL
XFILL_11_MUX2X1_24 gnd vdd FILL
XFILL_7_DFFSR_137 gnd vdd FILL
XDFFSR_151 DFFSR_151/Q CLKBUF1_6/Y DFFSR_23/R vdd DFFSR_151/D gnd vdd DFFSR
XFILL_11_MUX2X1_35 gnd vdd FILL
XBUFX4_3 rst_n gnd BUFX4_3/Y vdd BUFX4
XDFFSR_162 INVX1_147/A DFFSR_94/CLK DFFSR_99/R vdd MUX2X1_90/Y gnd vdd DFFSR
XFILL_7_DFFSR_148 gnd vdd FILL
XFILL_11_MUX2X1_46 gnd vdd FILL
XDFFSR_173 INVX1_90/A CLKBUF1_34/Y DFFSR_64/R vdd MUX2X1_35/Y gnd vdd DFFSR
XFILL_7_DFFSR_159 gnd vdd FILL
XFILL_11_MUX2X1_57 gnd vdd FILL
XDFFSR_184 INVX1_144/A DFFSR_99/CLK DFFSR_98/R vdd MUX2X1_1/Y gnd vdd DFFSR
XFILL_4_BUFX4_80 gnd vdd FILL
XFILL_4_BUFX4_91 gnd vdd FILL
XFILL_10_NOR3X1_9 gnd vdd FILL
XFILL_11_MUX2X1_68 gnd vdd FILL
XFILL_11_MUX2X1_79 gnd vdd FILL
XDFFSR_195 DFFSR_196/D CLKBUF1_7/Y BUFX4_13/Y vdd prev gnd vdd DFFSR
XFILL_15_MUX2X1_12 gnd vdd FILL
XFILL_15_MUX2X1_23 gnd vdd FILL
XFILL_41_DFFSR_190 gnd vdd FILL
XFILL_15_MUX2X1_34 gnd vdd FILL
XFILL_15_MUX2X1_45 gnd vdd FILL
XFILL_15_MUX2X1_56 gnd vdd FILL
XFILL_15_MUX2X1_67 gnd vdd FILL
XFILL_3_NOR3X1_16 gnd vdd FILL
XFILL_15_MUX2X1_78 gnd vdd FILL
XFILL_22_MUX2X1_1 gnd vdd FILL
XFILL_3_NOR3X1_27 gnd vdd FILL
XFILL_15_MUX2X1_89 gnd vdd FILL
XFILL_3_NOR3X1_38 gnd vdd FILL
XFILL_19_MUX2X1_11 gnd vdd FILL
XFILL_19_MUX2X1_22 gnd vdd FILL
XFILL_23_CLKBUF1_19 gnd vdd FILL
XFILL_3_NOR3X1_49 gnd vdd FILL
XFILL_19_MUX2X1_33 gnd vdd FILL
XFILL_19_MUX2X1_44 gnd vdd FILL
XFILL_57_4_0 gnd vdd FILL
XFILL_19_MUX2X1_55 gnd vdd FILL
XFILL_6_NOR2X1_4 gnd vdd FILL
XFILL_19_MUX2X1_66 gnd vdd FILL
XFILL_29_1_2 gnd vdd FILL
XFILL_19_MUX2X1_77 gnd vdd FILL
XFILL_4_1_2 gnd vdd FILL
XFILL_7_NOR3X1_15 gnd vdd FILL
XFILL_19_MUX2X1_88 gnd vdd FILL
XFILL_7_NOR3X1_26 gnd vdd FILL
XNOR3X1_40 NOR3X1_40/A NOR3X1_49/B NOR3X1_1/B gnd NOR3X1_42/A vdd NOR3X1
XFILL_19_MUX2X1_99 gnd vdd FILL
XNOR3X1_51 NOR3X1_9/A NOR3X1_9/B NOR3X1_51/C gnd NOR3X1_51/Y vdd NOR3X1
XFILL_8_MUX2X1_190 gnd vdd FILL
XFILL_7_NOR3X1_37 gnd vdd FILL
XFILL_23_DFFSR_102 gnd vdd FILL
XFILL_0_INVX1_109 gnd vdd FILL
XFILL_7_NOR3X1_48 gnd vdd FILL
XFILL_23_DFFSR_113 gnd vdd FILL
XFILL_23_DFFSR_124 gnd vdd FILL
XFILL_23_DFFSR_135 gnd vdd FILL
XFILL_23_DFFSR_146 gnd vdd FILL
XFILL_23_DFFSR_157 gnd vdd FILL
XFILL_23_DFFSR_168 gnd vdd FILL
XFILL_23_DFFSR_179 gnd vdd FILL
XFILL_5_MUX2X1_2 gnd vdd FILL
XFILL_4_INVX1_108 gnd vdd FILL
XFILL_27_DFFSR_101 gnd vdd FILL
XFILL_27_DFFSR_112 gnd vdd FILL
XFILL_4_INVX1_119 gnd vdd FILL
XFILL_4_NOR2X1_108 gnd vdd FILL
XFILL_27_DFFSR_123 gnd vdd FILL
XFILL_4_NOR2X1_119 gnd vdd FILL
XFILL_27_DFFSR_134 gnd vdd FILL
XFILL_31_DFFSR_4 gnd vdd FILL
XFILL_40_3_0 gnd vdd FILL
XFILL_27_DFFSR_145 gnd vdd FILL
XFILL_12_0_2 gnd vdd FILL
XFILL_10_NAND3X1_10 gnd vdd FILL
XFILL_27_DFFSR_156 gnd vdd FILL
XFILL_10_NAND3X1_21 gnd vdd FILL
XFILL_27_DFFSR_167 gnd vdd FILL
XFILL_10_NAND3X1_32 gnd vdd FILL
XFILL_27_DFFSR_178 gnd vdd FILL
XFILL_69_DFFSR_2 gnd vdd FILL
XFILL_10_NAND3X1_43 gnd vdd FILL
XFILL_27_DFFSR_189 gnd vdd FILL
XFILL_10_NAND3X1_54 gnd vdd FILL
XFILL_10_NAND3X1_65 gnd vdd FILL
XFILL_30_CLKBUF1_10 gnd vdd FILL
XFILL_30_CLKBUF1_21 gnd vdd FILL
XFILL_10_NAND3X1_76 gnd vdd FILL
XFILL_2_NOR3X1_8 gnd vdd FILL
XFILL_10_NAND3X1_87 gnd vdd FILL
XFILL_30_CLKBUF1_32 gnd vdd FILL
XFILL_10_NAND3X1_98 gnd vdd FILL
XFILL_39_DFFSR_80 gnd vdd FILL
XFILL_23_NOR3X1_13 gnd vdd FILL
XFILL_23_NOR3X1_24 gnd vdd FILL
XFILL_39_DFFSR_91 gnd vdd FILL
XFILL_23_NOR3X1_35 gnd vdd FILL
XFILL_23_NOR3X1_46 gnd vdd FILL
XFILL_73_DFFSR_202 gnd vdd FILL
XFILL_73_DFFSR_213 gnd vdd FILL
XFILL_0_DFFSR_10 gnd vdd FILL
XFILL_73_DFFSR_224 gnd vdd FILL
XFILL_73_DFFSR_235 gnd vdd FILL
XFILL_0_DFFSR_21 gnd vdd FILL
XFILL_0_DFFSR_32 gnd vdd FILL
XFILL_0_DFFSR_43 gnd vdd FILL
XFILL_73_DFFSR_246 gnd vdd FILL
XFILL_79_DFFSR_90 gnd vdd FILL
XFILL_27_NOR3X1_12 gnd vdd FILL
XFILL_0_DFFSR_54 gnd vdd FILL
XFILL_73_DFFSR_257 gnd vdd FILL
XFILL_73_DFFSR_268 gnd vdd FILL
XFILL_0_DFFSR_65 gnd vdd FILL
XFILL_27_NOR3X1_23 gnd vdd FILL
XFILL_27_NOR3X1_34 gnd vdd FILL
XFILL_53_DFFSR_8 gnd vdd FILL
XFILL_0_DFFSR_76 gnd vdd FILL
XFILL_27_NOR3X1_45 gnd vdd FILL
XFILL_77_DFFSR_201 gnd vdd FILL
XFILL_0_DFFSR_87 gnd vdd FILL
XFILL_0_DFFSR_98 gnd vdd FILL
XFILL_77_DFFSR_212 gnd vdd FILL
XFILL_77_DFFSR_223 gnd vdd FILL
XFILL_77_DFFSR_234 gnd vdd FILL
XFILL_1_OAI22X1_17 gnd vdd FILL
XFILL_77_DFFSR_245 gnd vdd FILL
XFILL_1_OAI22X1_28 gnd vdd FILL
XFILL_63_8 gnd vdd FILL
XFILL_77_DFFSR_256 gnd vdd FILL
XFILL_1_OAI22X1_39 gnd vdd FILL
XFILL_48_4_0 gnd vdd FILL
XFILL_77_DFFSR_267 gnd vdd FILL
XFILL_32_CLKBUF1_8 gnd vdd FILL
XFILL_14_AOI22X1_10 gnd vdd FILL
XFILL_5_OAI21X1_19 gnd vdd FILL
XFILL_0_NAND3X1_60 gnd vdd FILL
XFILL_0_NAND3X1_71 gnd vdd FILL
XFILL_0_NAND3X1_82 gnd vdd FILL
XFILL_4_NAND2X1_40 gnd vdd FILL
XFILL_0_NAND3X1_93 gnd vdd FILL
XFILL_4_NAND2X1_51 gnd vdd FILL
XFILL_4_NAND2X1_62 gnd vdd FILL
XFILL_4_NAND2X1_73 gnd vdd FILL
XFILL_4_NAND2X1_84 gnd vdd FILL
XFILL_4_NAND2X1_95 gnd vdd FILL
XFILL_31_3_0 gnd vdd FILL
XFILL_12_CLKBUF1_15 gnd vdd FILL
XFILL_12_CLKBUF1_26 gnd vdd FILL
XFILL_12_CLKBUF1_37 gnd vdd FILL
XFILL_10_NOR2X1_100 gnd vdd FILL
XFILL_10_NOR2X1_111 gnd vdd FILL
XFILL_10_NOR2X1_122 gnd vdd FILL
XFILL_10_NOR2X1_133 gnd vdd FILL
XFILL_10_NOR2X1_144 gnd vdd FILL
XFILL_10_NOR2X1_155 gnd vdd FILL
XFILL_10_NOR2X1_166 gnd vdd FILL
XFILL_40_DFFSR_202 gnd vdd FILL
XFILL_10_NOR2X1_177 gnd vdd FILL
XFILL_40_DFFSR_213 gnd vdd FILL
XFILL_10_NOR2X1_188 gnd vdd FILL
XFILL_2_OAI21X1_3 gnd vdd FILL
XFILL_10_NOR2X1_199 gnd vdd FILL
XFILL_40_DFFSR_224 gnd vdd FILL
XFILL_40_DFFSR_235 gnd vdd FILL
XFILL_8_AOI21X1_40 gnd vdd FILL
XFILL_40_DFFSR_246 gnd vdd FILL
XFILL_8_AOI21X1_51 gnd vdd FILL
XFILL_40_DFFSR_257 gnd vdd FILL
XFILL_40_DFFSR_268 gnd vdd FILL
XNAND3X1_6 DFFSR_22/Q BUFX4_8/Y NOR2X1_34/Y gnd NAND3X1_8/C vdd NAND3X1
XFILL_18_OAI22X1_20 gnd vdd FILL
XFILL_8_AOI21X1_62 gnd vdd FILL
XFILL_8_AOI21X1_73 gnd vdd FILL
XFILL_18_OAI22X1_31 gnd vdd FILL
XFILL_44_DFFSR_201 gnd vdd FILL
XFILL_18_OAI22X1_42 gnd vdd FILL
XFILL_44_DFFSR_212 gnd vdd FILL
XFILL_6_OAI21X1_2 gnd vdd FILL
XFILL_39_4_0 gnd vdd FILL
XFILL_44_DFFSR_223 gnd vdd FILL
XFILL_44_DFFSR_234 gnd vdd FILL
XFILL_3_NOR2X1_60 gnd vdd FILL
XFILL_44_DFFSR_245 gnd vdd FILL
XFILL_3_NOR2X1_71 gnd vdd FILL
XFILL_13_BUFX4_15 gnd vdd FILL
XFILL_2_CLKBUF1_10 gnd vdd FILL
XFILL_44_DFFSR_256 gnd vdd FILL
XFILL_2_CLKBUF1_21 gnd vdd FILL
XFILL_44_DFFSR_267 gnd vdd FILL
XFILL_3_NOR2X1_82 gnd vdd FILL
XFILL_2_CLKBUF1_32 gnd vdd FILL
XFILL_13_BUFX4_26 gnd vdd FILL
XFILL_71_DFFSR_101 gnd vdd FILL
XFILL_3_NOR2X1_93 gnd vdd FILL
XFILL_13_BUFX4_37 gnd vdd FILL
XFILL_48_DFFSR_200 gnd vdd FILL
XFILL_10_MUX2X1_106 gnd vdd FILL
XFILL_13_BUFX4_48 gnd vdd FILL
XFILL_71_DFFSR_112 gnd vdd FILL
XFILL_10_MUX2X1_117 gnd vdd FILL
XFILL_48_DFFSR_211 gnd vdd FILL
XFILL_13_BUFX4_59 gnd vdd FILL
XFILL_48_DFFSR_222 gnd vdd FILL
XFILL_71_DFFSR_123 gnd vdd FILL
XFILL_71_DFFSR_134 gnd vdd FILL
XFILL_48_DFFSR_233 gnd vdd FILL
XFILL_10_MUX2X1_128 gnd vdd FILL
XFILL_71_DFFSR_145 gnd vdd FILL
XFILL_10_MUX2X1_139 gnd vdd FILL
XFILL_48_DFFSR_244 gnd vdd FILL
XFILL_71_DFFSR_156 gnd vdd FILL
XFILL_48_DFFSR_255 gnd vdd FILL
XFILL_71_DFFSR_167 gnd vdd FILL
XFILL_7_NOR2X1_70 gnd vdd FILL
XFILL_7_NOR2X1_81 gnd vdd FILL
XFILL_48_DFFSR_266 gnd vdd FILL
XFILL_71_DFFSR_178 gnd vdd FILL
XFILL_7_NOR2X1_92 gnd vdd FILL
XFILL_75_DFFSR_100 gnd vdd FILL
XFILL_71_DFFSR_189 gnd vdd FILL
XFILL_75_DFFSR_111 gnd vdd FILL
XFILL_11_OAI21X1_11 gnd vdd FILL
XFILL_75_DFFSR_122 gnd vdd FILL
XFILL_11_OAI21X1_22 gnd vdd FILL
XFILL_0_DFFSR_3 gnd vdd FILL
XFILL_75_DFFSR_133 gnd vdd FILL
XFILL_11_OAI21X1_33 gnd vdd FILL
XFILL_22_3_0 gnd vdd FILL
XFILL_75_DFFSR_144 gnd vdd FILL
XFILL_11_OAI21X1_44 gnd vdd FILL
XFILL_75_DFFSR_155 gnd vdd FILL
XFILL_0_NOR2X1_150 gnd vdd FILL
XFILL_13_DFFSR_1 gnd vdd FILL
XFILL_0_NOR2X1_161 gnd vdd FILL
XFILL_75_DFFSR_166 gnd vdd FILL
XFILL_75_DFFSR_177 gnd vdd FILL
XFILL_70_DFFSR_2 gnd vdd FILL
XFILL_0_NOR2X1_172 gnd vdd FILL
XFILL_0_NOR2X1_183 gnd vdd FILL
XFILL_75_DFFSR_188 gnd vdd FILL
XFILL_0_NOR2X1_194 gnd vdd FILL
XFILL_79_DFFSR_110 gnd vdd FILL
XFILL_75_DFFSR_199 gnd vdd FILL
XFILL_79_DFFSR_121 gnd vdd FILL
XFILL_79_DFFSR_132 gnd vdd FILL
XFILL_79_DFFSR_143 gnd vdd FILL
XFILL_79_DFFSR_154 gnd vdd FILL
XFILL_7_INVX1_16 gnd vdd FILL
XFILL_79_DFFSR_165 gnd vdd FILL
XFILL_7_INVX1_27 gnd vdd FILL
XFILL_7_INVX1_38 gnd vdd FILL
XFILL_79_DFFSR_176 gnd vdd FILL
XFILL_79_DFFSR_187 gnd vdd FILL
XFILL_8_AND2X2_8 gnd vdd FILL
XFILL_7_INVX1_49 gnd vdd FILL
XFILL_79_DFFSR_198 gnd vdd FILL
XFILL_0_MUX2X1_101 gnd vdd FILL
XFILL_0_MUX2X1_112 gnd vdd FILL
XFILL_3_NAND2X1_4 gnd vdd FILL
XFILL_0_MUX2X1_123 gnd vdd FILL
XFILL_0_MUX2X1_134 gnd vdd FILL
XFILL_35_DFFSR_5 gnd vdd FILL
XFILL_0_MUX2X1_145 gnd vdd FILL
XFILL_5_BUFX4_14 gnd vdd FILL
XFILL_0_MUX2X1_156 gnd vdd FILL
XFILL_5_BUFX4_25 gnd vdd FILL
XFILL_0_MUX2X1_167 gnd vdd FILL
XFILL_5_BUFX4_36 gnd vdd FILL
XFILL_0_MUX2X1_178 gnd vdd FILL
XFILL_0_MUX2X1_189 gnd vdd FILL
XFILL_5_BUFX4_47 gnd vdd FILL
XFILL_5_BUFX4_58 gnd vdd FILL
XFILL_5_BUFX4_69 gnd vdd FILL
XFILL_5_4_0 gnd vdd FILL
XFILL_7_NAND2X1_3 gnd vdd FILL
XFILL_11_DFFSR_201 gnd vdd FILL
XFILL_11_DFFSR_212 gnd vdd FILL
XFILL_1_OAI21X1_50 gnd vdd FILL
XFILL_11_DFFSR_223 gnd vdd FILL
XFILL_11_DFFSR_234 gnd vdd FILL
XFILL_11_DFFSR_245 gnd vdd FILL
XFILL_11_DFFSR_256 gnd vdd FILL
XFILL_11_DFFSR_267 gnd vdd FILL
XFILL_15_DFFSR_200 gnd vdd FILL
XFILL_15_DFFSR_211 gnd vdd FILL
XFILL_15_DFFSR_222 gnd vdd FILL
XFILL_15_DFFSR_233 gnd vdd FILL
XFILL_15_DFFSR_244 gnd vdd FILL
XFILL_15_DFFSR_255 gnd vdd FILL
XFILL_15_DFFSR_266 gnd vdd FILL
XFILL_57_DFFSR_9 gnd vdd FILL
XFILL_13_3_0 gnd vdd FILL
XFILL_42_DFFSR_100 gnd vdd FILL
XFILL_42_DFFSR_111 gnd vdd FILL
XFILL_12_AND2X2_2 gnd vdd FILL
XFILL_19_DFFSR_210 gnd vdd FILL
XFILL_19_DFFSR_221 gnd vdd FILL
XFILL_42_DFFSR_122 gnd vdd FILL
XFILL_3_AOI21X1_9 gnd vdd FILL
XFILL_42_DFFSR_133 gnd vdd FILL
XFILL_19_DFFSR_232 gnd vdd FILL
XFILL_19_DFFSR_243 gnd vdd FILL
XFILL_42_DFFSR_144 gnd vdd FILL
XFILL_42_DFFSR_155 gnd vdd FILL
XFILL_19_DFFSR_254 gnd vdd FILL
XFILL_42_DFFSR_166 gnd vdd FILL
XFILL_19_DFFSR_265 gnd vdd FILL
XFILL_42_DFFSR_177 gnd vdd FILL
XFILL_42_DFFSR_188 gnd vdd FILL
XFILL_46_DFFSR_110 gnd vdd FILL
XFILL_42_DFFSR_199 gnd vdd FILL
XFILL_46_DFFSR_121 gnd vdd FILL
XFILL_3_NAND3X1_15 gnd vdd FILL
XFILL_46_DFFSR_132 gnd vdd FILL
XFILL_7_AOI21X1_8 gnd vdd FILL
XFILL_3_NAND3X1_26 gnd vdd FILL
XFILL_46_DFFSR_143 gnd vdd FILL
XFILL_3_NAND3X1_37 gnd vdd FILL
XFILL_46_DFFSR_154 gnd vdd FILL
XNOR3X1_9 NOR3X1_9/A NOR3X1_9/B NOR3X1_9/C gnd NOR3X1_9/Y vdd NOR3X1
XFILL_3_NAND3X1_48 gnd vdd FILL
XFILL_3_NAND3X1_59 gnd vdd FILL
XFILL_46_DFFSR_165 gnd vdd FILL
XFILL_46_DFFSR_176 gnd vdd FILL
XFILL_7_NAND2X1_17 gnd vdd FILL
XFILL_7_NAND2X1_28 gnd vdd FILL
XFILL_46_DFFSR_187 gnd vdd FILL
XFILL_7_NAND2X1_39 gnd vdd FILL
XFILL_46_DFFSR_198 gnd vdd FILL
XFILL_12_AOI22X1_5 gnd vdd FILL
XMUX2X1_180 BUFX4_66/Y OAI22X1_9/C NOR2X1_167/Y gnd DFFSR_60/D vdd MUX2X1
XMUX2X1_191 BUFX4_93/Y INVX1_11/Y NOR2X1_169/Y gnd DFFSR_53/D vdd MUX2X1
XFILL_5_3 gnd vdd FILL
XFILL_17_MUX2X1_170 gnd vdd FILL
XFILL_17_MUX2X1_181 gnd vdd FILL
XFILL_17_MUX2X1_192 gnd vdd FILL
XFILL_61_5 gnd vdd FILL
XFILL_16_AOI22X1_4 gnd vdd FILL
XFILL_54_4 gnd vdd FILL
XFILL_64_7_1 gnd vdd FILL
XFILL_11_NOR2X1_9 gnd vdd FILL
XFILL_63_2_0 gnd vdd FILL
XFILL_3_INVX1_20 gnd vdd FILL
XFILL_3_INVX1_31 gnd vdd FILL
XFILL_3_INVX1_42 gnd vdd FILL
XFILL_4_AND2X2_1 gnd vdd FILL
XFILL_3_INVX1_53 gnd vdd FILL
XFILL_3_INVX1_64 gnd vdd FILL
XFILL_49_DFFSR_12 gnd vdd FILL
XFILL_3_INVX1_75 gnd vdd FILL
XFILL_3_INVX1_86 gnd vdd FILL
XFILL_49_DFFSR_23 gnd vdd FILL
XFILL_3_INVX1_97 gnd vdd FILL
XFILL_49_DFFSR_34 gnd vdd FILL
XFILL_49_DFFSR_45 gnd vdd FILL
XFILL_49_DFFSR_56 gnd vdd FILL
XFILL_49_DFFSR_67 gnd vdd FILL
XFILL_10_MUX2X1_7 gnd vdd FILL
XFILL_49_DFFSR_78 gnd vdd FILL
XFILL_49_DFFSR_89 gnd vdd FILL
XFILL_22_CLKBUF1_16 gnd vdd FILL
XFILL_22_CLKBUF1_27 gnd vdd FILL
XFILL_22_CLKBUF1_38 gnd vdd FILL
XFILL_1_BUFX4_40 gnd vdd FILL
XFILL_1_BUFX4_51 gnd vdd FILL
XFILL_18_DFFSR_11 gnd vdd FILL
XFILL_18_DFFSR_22 gnd vdd FILL
XFILL_18_DFFSR_33 gnd vdd FILL
XFILL_1_BUFX4_62 gnd vdd FILL
XFILL_1_BUFX4_73 gnd vdd FILL
XFILL_18_DFFSR_44 gnd vdd FILL
XFILL_1_BUFX4_84 gnd vdd FILL
XFILL_1_BUFX4_95 gnd vdd FILL
XFILL_18_DFFSR_55 gnd vdd FILL
XFILL_18_DFFSR_66 gnd vdd FILL
XFILL_13_DFFSR_110 gnd vdd FILL
XFILL_18_DFFSR_77 gnd vdd FILL
XFILL_13_DFFSR_121 gnd vdd FILL
XFILL_0_AOI21X1_17 gnd vdd FILL
XFILL_18_DFFSR_88 gnd vdd FILL
XFILL_13_DFFSR_132 gnd vdd FILL
XFILL_18_DFFSR_99 gnd vdd FILL
XFILL_0_AOI21X1_28 gnd vdd FILL
XFILL_13_DFFSR_143 gnd vdd FILL
XFILL_0_AOI21X1_39 gnd vdd FILL
XFILL_58_DFFSR_10 gnd vdd FILL
XFILL_13_DFFSR_154 gnd vdd FILL
XFILL_58_DFFSR_21 gnd vdd FILL
XFILL_13_DFFSR_165 gnd vdd FILL
XFILL_58_DFFSR_32 gnd vdd FILL
XFILL_58_DFFSR_43 gnd vdd FILL
XFILL_10_OAI22X1_19 gnd vdd FILL
XFILL_29_NOR3X1_7 gnd vdd FILL
XFILL_2_CLKBUF1_8 gnd vdd FILL
XFILL_58_DFFSR_54 gnd vdd FILL
XFILL_13_DFFSR_176 gnd vdd FILL
XFILL_13_DFFSR_187 gnd vdd FILL
XFILL_13_DFFSR_198 gnd vdd FILL
XFILL_58_DFFSR_65 gnd vdd FILL
XFILL_58_DFFSR_76 gnd vdd FILL
XFILL_3_NOR2X1_105 gnd vdd FILL
XFILL_17_DFFSR_120 gnd vdd FILL
XFILL_17_DFFSR_131 gnd vdd FILL
XFILL_58_DFFSR_87 gnd vdd FILL
XFILL_3_NOR2X1_116 gnd vdd FILL
XFILL_4_DFFSR_4 gnd vdd FILL
XFILL_58_DFFSR_98 gnd vdd FILL
XFILL_3_NOR2X1_127 gnd vdd FILL
XFILL_17_DFFSR_142 gnd vdd FILL
XFILL_17_DFFSR_153 gnd vdd FILL
XFILL_17_DFFSR_2 gnd vdd FILL
XFILL_3_NOR2X1_138 gnd vdd FILL
XFILL_3_NOR2X1_149 gnd vdd FILL
XFILL_17_DFFSR_164 gnd vdd FILL
XFILL_17_DFFSR_175 gnd vdd FILL
XFILL_3_NOR2X1_8 gnd vdd FILL
XFILL_74_DFFSR_3 gnd vdd FILL
XFILL_6_CLKBUF1_7 gnd vdd FILL
XFILL_17_DFFSR_186 gnd vdd FILL
XFILL_17_DFFSR_197 gnd vdd FILL
XFILL_27_DFFSR_20 gnd vdd FILL
XFILL_27_DFFSR_31 gnd vdd FILL
XFILL_27_DFFSR_42 gnd vdd FILL
XFILL_27_DFFSR_53 gnd vdd FILL
XFILL_27_DFFSR_64 gnd vdd FILL
XFILL_2_BUFX4_102 gnd vdd FILL
XFILL_27_DFFSR_75 gnd vdd FILL
XFILL_55_7_1 gnd vdd FILL
XFILL_27_DFFSR_86 gnd vdd FILL
XFILL_13_NOR3X1_10 gnd vdd FILL
XFILL_27_DFFSR_97 gnd vdd FILL
XFILL_13_NOR3X1_21 gnd vdd FILL
XFILL_54_2_0 gnd vdd FILL
XFILL_13_NOR3X1_32 gnd vdd FILL
XFILL_67_DFFSR_30 gnd vdd FILL
XFILL_13_NOR3X1_43 gnd vdd FILL
XFILL_67_DFFSR_41 gnd vdd FILL
XFILL_2_MUX2X1_6 gnd vdd FILL
XFILL_20_MUX2X1_107 gnd vdd FILL
XFILL_63_DFFSR_210 gnd vdd FILL
XFILL_20_MUX2X1_118 gnd vdd FILL
XFILL_67_DFFSR_52 gnd vdd FILL
XFILL_67_DFFSR_63 gnd vdd FILL
XFILL_63_DFFSR_221 gnd vdd FILL
XFILL_20_MUX2X1_129 gnd vdd FILL
XFILL_6_BUFX4_101 gnd vdd FILL
XFILL_67_DFFSR_74 gnd vdd FILL
XFILL_63_DFFSR_232 gnd vdd FILL
XFILL_63_DFFSR_243 gnd vdd FILL
XFILL_67_DFFSR_85 gnd vdd FILL
XFILL_63_DFFSR_254 gnd vdd FILL
XFILL_67_DFFSR_96 gnd vdd FILL
XFILL_63_DFFSR_265 gnd vdd FILL
XFILL_17_NOR3X1_20 gnd vdd FILL
XFILL_17_NOR3X1_31 gnd vdd FILL
XFILL_17_NOR3X1_42 gnd vdd FILL
XFILL_39_DFFSR_6 gnd vdd FILL
XFILL_8_NOR2X1_205 gnd vdd FILL
XFILL_67_DFFSR_220 gnd vdd FILL
XFILL_0_OAI22X1_14 gnd vdd FILL
XFILL_67_DFFSR_231 gnd vdd FILL
XFILL_67_DFFSR_242 gnd vdd FILL
XFILL_0_OAI22X1_25 gnd vdd FILL
XFILL_36_DFFSR_40 gnd vdd FILL
XFILL_0_OAI22X1_36 gnd vdd FILL
XFILL_36_DFFSR_51 gnd vdd FILL
XFILL_67_DFFSR_253 gnd vdd FILL
XFILL_0_OAI22X1_47 gnd vdd FILL
XFILL_36_DFFSR_62 gnd vdd FILL
XFILL_67_DFFSR_264 gnd vdd FILL
XFILL_67_DFFSR_275 gnd vdd FILL
XFILL_4_OAI21X1_16 gnd vdd FILL
XFILL_36_DFFSR_73 gnd vdd FILL
XFILL_22_CLKBUF1_5 gnd vdd FILL
XFILL_36_DFFSR_84 gnd vdd FILL
XFILL_4_OAI21X1_27 gnd vdd FILL
XFILL_0_NOR2X1_15 gnd vdd FILL
XFILL_0_NOR2X1_26 gnd vdd FILL
XFILL_36_DFFSR_95 gnd vdd FILL
XAOI21X1_30 BUFX4_83/Y NOR2X1_190/B NOR2X1_187/Y gnd DFFSR_19/D vdd AOI21X1
XFILL_4_OAI21X1_38 gnd vdd FILL
XFILL_4_OAI21X1_49 gnd vdd FILL
XAOI21X1_41 BUFX4_71/Y NOR2X1_202/B NOR2X1_201/Y gnd DFFSR_8/D vdd AOI21X1
XFILL_0_NOR2X1_37 gnd vdd FILL
XAOI21X1_52 MUX2X1_8/A NOR2X1_12/B NOR2X1_11/Y gnd DFFSR_262/D vdd AOI21X1
XFILL_0_NOR2X1_48 gnd vdd FILL
XFILL_0_NOR2X1_59 gnd vdd FILL
XAOI21X1_63 OAI21X1_45/Y NAND3X1_39/B NAND3X1_43/A gnd AND2X2_5/B vdd AOI21X1
XAOI21X1_74 INVX1_104/A INVX1_125/Y OAI22X1_41/Y gnd NAND3X1_18/B vdd AOI21X1
XFILL_76_DFFSR_50 gnd vdd FILL
XFILL_26_CLKBUF1_4 gnd vdd FILL
XFILL_76_DFFSR_61 gnd vdd FILL
XFILL_76_DFFSR_72 gnd vdd FILL
XFILL_76_DFFSR_83 gnd vdd FILL
XOAI21X1_3 OAI21X1_3/A OAI21X1_3/B OAI21X1_3/C gnd OAI21X1_3/Y vdd OAI21X1
XFILL_76_DFFSR_94 gnd vdd FILL
XFILL_4_NOR2X1_14 gnd vdd FILL
XFILL_4_NOR2X1_25 gnd vdd FILL
XFILL_11_BUFX4_2 gnd vdd FILL
XFILL_3_NAND2X1_70 gnd vdd FILL
XFILL_3_NAND2X1_81 gnd vdd FILL
XFILL_4_NOR2X1_36 gnd vdd FILL
XFILL_4_NOR2X1_47 gnd vdd FILL
XFILL_3_NAND2X1_92 gnd vdd FILL
XFILL_4_NOR2X1_58 gnd vdd FILL
XFILL_9_0_2 gnd vdd FILL
XFILL_4_NOR2X1_69 gnd vdd FILL
XFILL_11_CLKBUF1_12 gnd vdd FILL
XFILL_16_NOR3X1_2 gnd vdd FILL
XFILL_11_CLKBUF1_23 gnd vdd FILL
XFILL_8_NOR2X1_13 gnd vdd FILL
XFILL_8_NOR2X1_24 gnd vdd FILL
XFILL_49_DFFSR_209 gnd vdd FILL
XFILL_11_CLKBUF1_34 gnd vdd FILL
XFILL_45_DFFSR_60 gnd vdd FILL
XFILL_8_NOR2X1_35 gnd vdd FILL
XFILL_45_DFFSR_71 gnd vdd FILL
XFILL_45_DFFSR_82 gnd vdd FILL
XFILL_8_NOR2X1_46 gnd vdd FILL
XFILL_12_OAI22X1_8 gnd vdd FILL
XFILL_45_DFFSR_93 gnd vdd FILL
XFILL_8_NOR2X1_57 gnd vdd FILL
XFILL_8_NOR2X1_68 gnd vdd FILL
XFILL_8_NOR2X1_79 gnd vdd FILL
XFILL_76_DFFSR_109 gnd vdd FILL
XFILL_46_7_1 gnd vdd FILL
XFILL_85_DFFSR_70 gnd vdd FILL
XFILL_45_2_0 gnd vdd FILL
XFILL_85_DFFSR_81 gnd vdd FILL
XFILL_85_DFFSR_92 gnd vdd FILL
XFILL_16_OAI22X1_7 gnd vdd FILL
XFILL_14_DFFSR_70 gnd vdd FILL
XFILL_14_DFFSR_81 gnd vdd FILL
XFILL_14_DFFSR_92 gnd vdd FILL
XFILL_30_DFFSR_210 gnd vdd FILL
XFILL_30_DFFSR_221 gnd vdd FILL
XFILL_26_8 gnd vdd FILL
XFILL_30_DFFSR_232 gnd vdd FILL
XFILL_30_DFFSR_243 gnd vdd FILL
XFILL_30_DFFSR_254 gnd vdd FILL
XFILL_30_DFFSR_265 gnd vdd FILL
XFILL_54_DFFSR_80 gnd vdd FILL
XFILL_7_AOI21X1_70 gnd vdd FILL
XFILL_7_AOI21X1_81 gnd vdd FILL
XFILL_54_DFFSR_91 gnd vdd FILL
XFILL_17_OAI22X1_50 gnd vdd FILL
XFILL_34_DFFSR_220 gnd vdd FILL
XFILL_34_DFFSR_231 gnd vdd FILL
XFILL_34_DFFSR_242 gnd vdd FILL
XFILL_34_DFFSR_253 gnd vdd FILL
XFILL_34_DFFSR_264 gnd vdd FILL
XFILL_0_MUX2X1_11 gnd vdd FILL
XFILL_34_DFFSR_275 gnd vdd FILL
XFILL_0_MUX2X1_22 gnd vdd FILL
XFILL_1_CLKBUF1_40 gnd vdd FILL
XFILL_1_INVX8_2 gnd vdd FILL
XFILL_0_MUX2X1_33 gnd vdd FILL
XFILL_61_DFFSR_120 gnd vdd FILL
XFILL_0_MUX2X1_44 gnd vdd FILL
XFILL_0_MUX2X1_55 gnd vdd FILL
XFILL_61_DFFSR_131 gnd vdd FILL
XFILL_0_MUX2X1_66 gnd vdd FILL
XFILL_38_DFFSR_230 gnd vdd FILL
XFILL_0_MUX2X1_77 gnd vdd FILL
XFILL_23_DFFSR_90 gnd vdd FILL
XFILL_61_DFFSR_142 gnd vdd FILL
XFILL_38_DFFSR_241 gnd vdd FILL
XFILL_61_DFFSR_153 gnd vdd FILL
XFILL_8_NOR3X1_1 gnd vdd FILL
XFILL_38_DFFSR_252 gnd vdd FILL
XFILL_0_MUX2X1_88 gnd vdd FILL
XFILL_61_DFFSR_164 gnd vdd FILL
XFILL_0_MUX2X1_99 gnd vdd FILL
XFILL_61_DFFSR_175 gnd vdd FILL
XFILL_4_MUX2X1_10 gnd vdd FILL
XFILL_38_DFFSR_263 gnd vdd FILL
XFILL_38_DFFSR_274 gnd vdd FILL
XFILL_4_MUX2X1_21 gnd vdd FILL
XFILL_61_DFFSR_186 gnd vdd FILL
XFILL_4_MUX2X1_32 gnd vdd FILL
XFILL_61_DFFSR_197 gnd vdd FILL
XFILL_4_MUX2X1_43 gnd vdd FILL
XFILL_65_DFFSR_130 gnd vdd FILL
XFILL_4_MUX2X1_54 gnd vdd FILL
XFILL_10_OAI21X1_30 gnd vdd FILL
XFILL_4_MUX2X1_65 gnd vdd FILL
XFILL_4_MUX2X1_76 gnd vdd FILL
XFILL_10_OAI21X1_41 gnd vdd FILL
XFILL_65_DFFSR_141 gnd vdd FILL
XFILL_65_DFFSR_152 gnd vdd FILL
XFILL_4_MUX2X1_87 gnd vdd FILL
XFILL_65_DFFSR_163 gnd vdd FILL
XFILL_65_DFFSR_174 gnd vdd FILL
XFILL_4_MUX2X1_98 gnd vdd FILL
XFILL_8_MUX2X1_20 gnd vdd FILL
XFILL_65_DFFSR_185 gnd vdd FILL
XFILL_8_MUX2X1_31 gnd vdd FILL
XFILL_8_MUX2X1_42 gnd vdd FILL
XFILL_10_BUFX4_19 gnd vdd FILL
XFILL_65_DFFSR_196 gnd vdd FILL
XFILL_13_NAND3X1_9 gnd vdd FILL
XFILL_16_DFFSR_209 gnd vdd FILL
XFILL_8_MUX2X1_53 gnd vdd FILL
XFILL_69_DFFSR_140 gnd vdd FILL
XFILL_8_MUX2X1_64 gnd vdd FILL
XFILL_6_DFFSR_80 gnd vdd FILL
XFILL_8_MUX2X1_75 gnd vdd FILL
XFILL_8_MUX2X1_86 gnd vdd FILL
XFILL_69_DFFSR_151 gnd vdd FILL
XFILL_69_DFFSR_162 gnd vdd FILL
XFILL_37_7_1 gnd vdd FILL
XFILL_6_DFFSR_91 gnd vdd FILL
XFILL_8_MUX2X1_97 gnd vdd FILL
XFILL_69_DFFSR_173 gnd vdd FILL
XFILL_69_DFFSR_184 gnd vdd FILL
XFILL_36_2_0 gnd vdd FILL
XFILL_43_DFFSR_109 gnd vdd FILL
XFILL_69_DFFSR_195 gnd vdd FILL
XFILL_47_DFFSR_108 gnd vdd FILL
XFILL_40_DFFSR_6 gnd vdd FILL
XFILL_47_DFFSR_119 gnd vdd FILL
XFILL_8_DFFSR_5 gnd vdd FILL
XFILL_20_MUX2X1_30 gnd vdd FILL
XFILL_20_MUX2X1_41 gnd vdd FILL
XFILL_20_MUX2X1_52 gnd vdd FILL
XFILL_12_NAND3X1_17 gnd vdd FILL
XFILL_20_MUX2X1_63 gnd vdd FILL
XFILL_12_NAND3X1_28 gnd vdd FILL
XFILL_20_MUX2X1_74 gnd vdd FILL
XFILL_78_DFFSR_4 gnd vdd FILL
XFILL_20_6_1 gnd vdd FILL
XFILL_12_NAND3X1_39 gnd vdd FILL
XFILL_20_MUX2X1_85 gnd vdd FILL
XFILL_20_MUX2X1_96 gnd vdd FILL
XFILL_32_CLKBUF1_17 gnd vdd FILL
XFILL_32_CLKBUF1_28 gnd vdd FILL
XFILL_32_CLKBUF1_39 gnd vdd FILL
XFILL_2_BUFX4_18 gnd vdd FILL
XFILL_2_BUFX4_29 gnd vdd FILL
XFILL_32_DFFSR_130 gnd vdd FILL
XFILL_32_DFFSR_141 gnd vdd FILL
XFILL_32_DFFSR_152 gnd vdd FILL
XFILL_32_DFFSR_163 gnd vdd FILL
XFILL_32_DFFSR_174 gnd vdd FILL
XFILL_32_DFFSR_185 gnd vdd FILL
XFILL_32_DFFSR_196 gnd vdd FILL
XFILL_2_NAND3X1_12 gnd vdd FILL
XFILL_3_7_1 gnd vdd FILL
XFILL_28_7_1 gnd vdd FILL
XFILL_2_NAND3X1_23 gnd vdd FILL
XFILL_36_DFFSR_140 gnd vdd FILL
XFILL_2_NAND3X1_34 gnd vdd FILL
XFILL_36_DFFSR_151 gnd vdd FILL
XFILL_2_2_0 gnd vdd FILL
XFILL_2_NAND3X1_45 gnd vdd FILL
XFILL_27_2_0 gnd vdd FILL
XFILL_36_DFFSR_162 gnd vdd FILL
XFILL_2_NAND3X1_56 gnd vdd FILL
XFILL_6_NAND2X1_14 gnd vdd FILL
XFILL_36_DFFSR_173 gnd vdd FILL
XFILL_2_NAND3X1_67 gnd vdd FILL
XFILL_36_DFFSR_184 gnd vdd FILL
XFILL_6_NAND2X1_25 gnd vdd FILL
XFILL_2_NAND3X1_78 gnd vdd FILL
XFILL_6_NAND2X1_36 gnd vdd FILL
XFILL_10_DFFSR_109 gnd vdd FILL
XFILL_2_NAND3X1_89 gnd vdd FILL
XFILL_36_DFFSR_195 gnd vdd FILL
XFILL_6_NAND2X1_47 gnd vdd FILL
XFILL_2_BUFX4_5 gnd vdd FILL
XFILL_15_BUFX4_3 gnd vdd FILL
XFILL_6_NAND2X1_58 gnd vdd FILL
XFILL_6_NAND2X1_69 gnd vdd FILL
XMUX2X1_7 MUX2X1_7/A MUX2X1_7/B MUX2X1_7/S gnd MUX2X1_7/Y vdd MUX2X1
XFILL_14_DFFSR_108 gnd vdd FILL
XFILL_14_DFFSR_119 gnd vdd FILL
XFILL_11_6_1 gnd vdd FILL
XFILL_68_DFFSR_19 gnd vdd FILL
XFILL_82_DFFSR_230 gnd vdd FILL
XFILL_10_1_0 gnd vdd FILL
XFILL_82_DFFSR_241 gnd vdd FILL
XFILL_82_DFFSR_252 gnd vdd FILL
XFILL_82_DFFSR_263 gnd vdd FILL
XFILL_82_DFFSR_274 gnd vdd FILL
XFILL_18_DFFSR_107 gnd vdd FILL
XFILL_18_DFFSR_118 gnd vdd FILL
XFILL_1_INVX1_9 gnd vdd FILL
XFILL_18_DFFSR_129 gnd vdd FILL
XFILL_13_AOI21X1_3 gnd vdd FILL
XCLKBUF1_8 BUFX4_84/Y gnd CLKBUF1_8/Y vdd CLKBUF1
XFILL_86_DFFSR_240 gnd vdd FILL
XFILL_86_DFFSR_251 gnd vdd FILL
XFILL_86_DFFSR_262 gnd vdd FILL
XFILL_37_DFFSR_18 gnd vdd FILL
XFILL_86_DFFSR_273 gnd vdd FILL
XFILL_37_DFFSR_29 gnd vdd FILL
XFILL_60_DFFSR_209 gnd vdd FILL
XFILL_2_INVX1_190 gnd vdd FILL
XFILL_77_DFFSR_17 gnd vdd FILL
XFILL_14_NOR3X1_19 gnd vdd FILL
XFILL_77_DFFSR_28 gnd vdd FILL
XFILL_21_CLKBUF1_13 gnd vdd FILL
XFILL_21_CLKBUF1_24 gnd vdd FILL
XFILL_77_DFFSR_39 gnd vdd FILL
XFILL_64_DFFSR_208 gnd vdd FILL
XFILL_21_CLKBUF1_35 gnd vdd FILL
XFILL_64_DFFSR_219 gnd vdd FILL
XBUFX4_102 BUFX4_2/A gnd BUFX4_102/Y vdd BUFX4
XFILL_0_INVX1_13 gnd vdd FILL
XFILL_19_7_1 gnd vdd FILL
XFILL_0_INVX1_24 gnd vdd FILL
XFILL_0_INVX1_35 gnd vdd FILL
XFILL_18_NOR3X1_18 gnd vdd FILL
XFILL_4_CLKBUF1_17 gnd vdd FILL
XFILL_4_CLKBUF1_28 gnd vdd FILL
XFILL_0_INVX1_46 gnd vdd FILL
XFILL_1_AND2X2_5 gnd vdd FILL
XFILL_18_NOR3X1_29 gnd vdd FILL
XFILL_18_2_0 gnd vdd FILL
XFILL_0_INVX1_57 gnd vdd FILL
XFILL_4_CLKBUF1_39 gnd vdd FILL
XFILL_5_INVX8_3 gnd vdd FILL
XNOR2X1_206 NOR2X1_27/A NOR2X1_7/B gnd NOR2X1_6/B vdd NOR2X1
XFILL_0_INVX1_68 gnd vdd FILL
XFILL_68_DFFSR_207 gnd vdd FILL
XFILL_18_INVX8_1 gnd vdd FILL
XFILL_46_DFFSR_16 gnd vdd FILL
XFILL_68_DFFSR_218 gnd vdd FILL
XFILL_0_INVX1_79 gnd vdd FILL
XFILL_46_DFFSR_27 gnd vdd FILL
XFILL_68_DFFSR_229 gnd vdd FILL
XFILL_46_DFFSR_38 gnd vdd FILL
XFILL_31_6 gnd vdd FILL
XFILL_61_5_1 gnd vdd FILL
XFILL_46_DFFSR_49 gnd vdd FILL
XFILL_60_0_0 gnd vdd FILL
XFILL_2_NOR2X1_102 gnd vdd FILL
XFILL_24_5 gnd vdd FILL
XFILL_2_NOR2X1_113 gnd vdd FILL
XFILL_2_NOR2X1_124 gnd vdd FILL
XFILL_13_OAI21X1_18 gnd vdd FILL
XFILL_86_DFFSR_15 gnd vdd FILL
XFILL_13_OAI21X1_29 gnd vdd FILL
XFILL_86_DFFSR_26 gnd vdd FILL
XFILL_2_NOR2X1_135 gnd vdd FILL
XFILL_22_DFFSR_3 gnd vdd FILL
XFILL_86_DFFSR_37 gnd vdd FILL
XFILL_17_4 gnd vdd FILL
XFILL_2_NOR2X1_146 gnd vdd FILL
XFILL_86_DFFSR_48 gnd vdd FILL
XFILL_2_NOR2X1_157 gnd vdd FILL
XFILL_15_DFFSR_15 gnd vdd FILL
XFILL_86_DFFSR_59 gnd vdd FILL
XFILL_2_NOR2X1_168 gnd vdd FILL
XFILL_15_DFFSR_26 gnd vdd FILL
XFILL_2_NOR2X1_179 gnd vdd FILL
XFILL_15_DFFSR_37 gnd vdd FILL
XFILL_15_DFFSR_48 gnd vdd FILL
XFILL_26_15 gnd vdd FILL
XFILL_15_DFFSR_59 gnd vdd FILL
XFILL_55_DFFSR_14 gnd vdd FILL
XFILL_55_DFFSR_25 gnd vdd FILL
XFILL_55_DFFSR_36 gnd vdd FILL
XFILL_55_DFFSR_47 gnd vdd FILL
XFILL_55_DFFSR_58 gnd vdd FILL
XFILL_55_DFFSR_69 gnd vdd FILL
XFILL_53_DFFSR_240 gnd vdd FILL
XFILL_53_DFFSR_251 gnd vdd FILL
XFILL_53_DFFSR_262 gnd vdd FILL
XFILL_53_DFFSR_273 gnd vdd FILL
XFILL_2_MUX2X1_108 gnd vdd FILL
XFILL_2_MUX2X1_119 gnd vdd FILL
XFILL_24_DFFSR_13 gnd vdd FILL
XFILL_44_DFFSR_7 gnd vdd FILL
XFILL_7_NOR2X1_202 gnd vdd FILL
XFILL_24_DFFSR_24 gnd vdd FILL
XFILL_24_DFFSR_35 gnd vdd FILL
XFILL_80_DFFSR_140 gnd vdd FILL
XFILL_24_DFFSR_46 gnd vdd FILL
XFILL_24_DFFSR_57 gnd vdd FILL
XFILL_80_DFFSR_151 gnd vdd FILL
XFILL_57_DFFSR_250 gnd vdd FILL
XFILL_80_DFFSR_162 gnd vdd FILL
XFILL_24_DFFSR_68 gnd vdd FILL
XFILL_80_DFFSR_173 gnd vdd FILL
XFILL_12_CLKBUF1_2 gnd vdd FILL
XFILL_57_DFFSR_261 gnd vdd FILL
XFILL_3_OAI21X1_13 gnd vdd FILL
XFILL_57_DFFSR_272 gnd vdd FILL
XFILL_24_DFFSR_79 gnd vdd FILL
XFILL_80_DFFSR_184 gnd vdd FILL
XFILL_3_OAI21X1_24 gnd vdd FILL
XFILL_0_DFFSR_210 gnd vdd FILL
XFILL_64_DFFSR_12 gnd vdd FILL
XFILL_80_DFFSR_195 gnd vdd FILL
XFILL_31_DFFSR_208 gnd vdd FILL
XFILL_3_OAI21X1_35 gnd vdd FILL
XFILL_0_DFFSR_221 gnd vdd FILL
XFILL_64_DFFSR_23 gnd vdd FILL
XFILL_31_DFFSR_219 gnd vdd FILL
XFILL_0_DFFSR_232 gnd vdd FILL
XFILL_3_OAI21X1_46 gnd vdd FILL
XFILL_0_DFFSR_243 gnd vdd FILL
XFILL_64_DFFSR_34 gnd vdd FILL
XFILL_64_DFFSR_45 gnd vdd FILL
XFILL_64_DFFSR_56 gnd vdd FILL
XFILL_0_DFFSR_254 gnd vdd FILL
XFILL_84_DFFSR_150 gnd vdd FILL
XFILL_84_DFFSR_161 gnd vdd FILL
XFILL_64_DFFSR_67 gnd vdd FILL
XFILL_0_DFFSR_265 gnd vdd FILL
XFILL_64_DFFSR_78 gnd vdd FILL
XFILL_16_CLKBUF1_1 gnd vdd FILL
XFILL_84_DFFSR_172 gnd vdd FILL
XFILL_84_DFFSR_183 gnd vdd FILL
XFILL_64_DFFSR_89 gnd vdd FILL
XFILL_84_DFFSR_194 gnd vdd FILL
XFILL_35_DFFSR_207 gnd vdd FILL
XFILL_4_DFFSR_220 gnd vdd FILL
XFILL_52_5_1 gnd vdd FILL
XFILL_7_DFFSR_14 gnd vdd FILL
XFILL_35_DFFSR_218 gnd vdd FILL
XFILL_4_DFFSR_231 gnd vdd FILL
XFILL_4_DFFSR_242 gnd vdd FILL
XFILL_35_DFFSR_229 gnd vdd FILL
XFILL_51_0_0 gnd vdd FILL
XFILL_7_DFFSR_25 gnd vdd FILL
XFILL_33_DFFSR_11 gnd vdd FILL
XFILL_7_DFFSR_36 gnd vdd FILL
XFILL_4_DFFSR_253 gnd vdd FILL
XFILL_33_DFFSR_22 gnd vdd FILL
XFILL_4_DFFSR_264 gnd vdd FILL
XFILL_7_DFFSR_47 gnd vdd FILL
XFILL_4_DFFSR_275 gnd vdd FILL
XFILL_7_DFFSR_58 gnd vdd FILL
XFILL_33_DFFSR_33 gnd vdd FILL
XFILL_7_DFFSR_69 gnd vdd FILL
XFILL_33_DFFSR_44 gnd vdd FILL
XFILL_39_DFFSR_206 gnd vdd FILL
XFILL_62_DFFSR_107 gnd vdd FILL
XFILL_10_CLKBUF1_20 gnd vdd FILL
XFILL_33_DFFSR_55 gnd vdd FILL
XFILL_33_DFFSR_66 gnd vdd FILL
XFILL_10_CLKBUF1_31 gnd vdd FILL
XFILL_62_DFFSR_118 gnd vdd FILL
XFILL_33_DFFSR_77 gnd vdd FILL
XFILL_39_DFFSR_217 gnd vdd FILL
XFILL_8_DFFSR_230 gnd vdd FILL
XFILL_8_DFFSR_241 gnd vdd FILL
XFILL_10_CLKBUF1_42 gnd vdd FILL
XFILL_39_DFFSR_228 gnd vdd FILL
XFILL_33_DFFSR_88 gnd vdd FILL
XFILL_62_DFFSR_129 gnd vdd FILL
XFILL_39_DFFSR_239 gnd vdd FILL
XFILL_8_DFFSR_252 gnd vdd FILL
XFILL_33_DFFSR_99 gnd vdd FILL
XFILL_73_DFFSR_10 gnd vdd FILL
XFILL_9_BUFX2_10 gnd vdd FILL
XFILL_73_DFFSR_21 gnd vdd FILL
XFILL_8_DFFSR_263 gnd vdd FILL
XFILL_8_DFFSR_274 gnd vdd FILL
XFILL_73_DFFSR_32 gnd vdd FILL
XFILL_73_DFFSR_43 gnd vdd FILL
XFILL_5_MUX2X1_19 gnd vdd FILL
XFILL_66_DFFSR_106 gnd vdd FILL
XFILL_73_DFFSR_54 gnd vdd FILL
XFILL_73_DFFSR_65 gnd vdd FILL
XFILL_66_DFFSR_117 gnd vdd FILL
XFILL_73_DFFSR_76 gnd vdd FILL
XFILL_66_DFFSR_128 gnd vdd FILL
XFILL_73_DFFSR_87 gnd vdd FILL
XFILL_73_DFFSR_98 gnd vdd FILL
XFILL_66_DFFSR_139 gnd vdd FILL
XFILL_9_MUX2X1_18 gnd vdd FILL
XFILL_9_MUX2X1_29 gnd vdd FILL
XFILL_6_BUFX4_6 gnd vdd FILL
XFILL_42_DFFSR_20 gnd vdd FILL
XFILL_19_MUX2X1_100 gnd vdd FILL
XFILL_42_DFFSR_31 gnd vdd FILL
XFILL_19_MUX2X1_111 gnd vdd FILL
XFILL_13_NOR3X1_6 gnd vdd FILL
XFILL_42_DFFSR_42 gnd vdd FILL
XFILL_10_NOR2X1_20 gnd vdd FILL
XFILL_19_MUX2X1_122 gnd vdd FILL
XFILL_10_NOR2X1_31 gnd vdd FILL
XFILL_42_DFFSR_53 gnd vdd FILL
XFILL_1_AOI22X1_3 gnd vdd FILL
XFILL_13_OAI21X1_6 gnd vdd FILL
XFILL_20_DFFSR_240 gnd vdd FILL
XFILL_19_MUX2X1_133 gnd vdd FILL
XFILL_10_NOR2X1_42 gnd vdd FILL
XFILL_42_DFFSR_64 gnd vdd FILL
XFILL_19_MUX2X1_144 gnd vdd FILL
XFILL_10_NOR2X1_53 gnd vdd FILL
XFILL_20_DFFSR_251 gnd vdd FILL
XFILL_42_DFFSR_75 gnd vdd FILL
XFILL_19_MUX2X1_155 gnd vdd FILL
XFILL_42_DFFSR_86 gnd vdd FILL
XFILL_20_DFFSR_262 gnd vdd FILL
XFILL_10_NOR2X1_64 gnd vdd FILL
XFILL_10_NOR2X1_75 gnd vdd FILL
XFILL_20_DFFSR_273 gnd vdd FILL
XFILL_19_MUX2X1_166 gnd vdd FILL
XFILL_42_DFFSR_97 gnd vdd FILL
XFILL_59_1_0 gnd vdd FILL
XFILL_1_INVX1_202 gnd vdd FILL
XBUFX4_19 BUFX4_62/Y gnd DFFSR_99/R vdd BUFX4
XFILL_19_MUX2X1_177 gnd vdd FILL
XFILL_19_MUX2X1_188 gnd vdd FILL
XFILL_1_INVX1_213 gnd vdd FILL
XFILL_10_NOR2X1_86 gnd vdd FILL
XFILL_82_DFFSR_30 gnd vdd FILL
XFILL_10_NOR2X1_97 gnd vdd FILL
XFILL_1_INVX1_224 gnd vdd FILL
XFILL_5_AOI22X1_2 gnd vdd FILL
XFILL_82_DFFSR_41 gnd vdd FILL
XFILL_82_DFFSR_52 gnd vdd FILL
XFILL_82_DFFSR_63 gnd vdd FILL
XFILL_24_DFFSR_250 gnd vdd FILL
XFILL_82_DFFSR_74 gnd vdd FILL
XFILL_11_DFFSR_30 gnd vdd FILL
XFILL_82_DFFSR_85 gnd vdd FILL
XFILL_11_DFFSR_41 gnd vdd FILL
XFILL_24_DFFSR_261 gnd vdd FILL
XFILL_24_DFFSR_272 gnd vdd FILL
XFILL_82_DFFSR_96 gnd vdd FILL
XFILL_11_DFFSR_52 gnd vdd FILL
XFILL_5_INVX1_201 gnd vdd FILL
XFILL_11_DFFSR_63 gnd vdd FILL
XFILL_21_MUX2X1_17 gnd vdd FILL
XFILL_5_INVX1_212 gnd vdd FILL
XFILL_9_NOR2X1_1 gnd vdd FILL
XFILL_21_MUX2X1_28 gnd vdd FILL
XFILL_5_INVX1_223 gnd vdd FILL
XFILL_11_DFFSR_74 gnd vdd FILL
XFILL_11_DFFSR_85 gnd vdd FILL
XFILL_21_MUX2X1_39 gnd vdd FILL
XFILL_9_AOI22X1_1 gnd vdd FILL
XFILL_11_DFFSR_96 gnd vdd FILL
XFILL_51_DFFSR_150 gnd vdd FILL
XFILL_51_DFFSR_161 gnd vdd FILL
XFILL_28_DFFSR_260 gnd vdd FILL
XFILL_51_DFFSR_40 gnd vdd FILL
XFILL_2_BUFX2_2 gnd vdd FILL
XFILL_43_5_1 gnd vdd FILL
XFILL_51_DFFSR_172 gnd vdd FILL
XFILL_22_NOR3X1_4 gnd vdd FILL
XFILL_28_DFFSR_271 gnd vdd FILL
XFILL_51_DFFSR_51 gnd vdd FILL
XFILL_51_DFFSR_183 gnd vdd FILL
XFILL_51_DFFSR_62 gnd vdd FILL
XFILL_42_0_0 gnd vdd FILL
XFILL_51_DFFSR_73 gnd vdd FILL
XFILL_51_DFFSR_194 gnd vdd FILL
XFILL_51_DFFSR_84 gnd vdd FILL
XFILL_51_DFFSR_95 gnd vdd FILL
XFILL_55_DFFSR_160 gnd vdd FILL
XFILL_55_DFFSR_171 gnd vdd FILL
XFILL_55_DFFSR_182 gnd vdd FILL
XFILL_61_DFFSR_1 gnd vdd FILL
XFILL_55_DFFSR_193 gnd vdd FILL
XFILL_20_DFFSR_50 gnd vdd FILL
XFILL_9_MUX2X1_150 gnd vdd FILL
XFILL_20_DFFSR_61 gnd vdd FILL
XFILL_9_MUX2X1_161 gnd vdd FILL
XFILL_20_DFFSR_72 gnd vdd FILL
XFILL_20_DFFSR_83 gnd vdd FILL
XFILL_59_DFFSR_170 gnd vdd FILL
XFILL_9_MUX2X1_172 gnd vdd FILL
XFILL_20_DFFSR_94 gnd vdd FILL
XFILL_9_MUX2X1_183 gnd vdd FILL
XFILL_59_DFFSR_181 gnd vdd FILL
XFILL_9_INVX8_4 gnd vdd FILL
XFILL_9_MUX2X1_194 gnd vdd FILL
XFILL_59_DFFSR_192 gnd vdd FILL
XFILL_5_NOR3X1_5 gnd vdd FILL
XFILL_33_DFFSR_106 gnd vdd FILL
XFILL_2_DFFSR_130 gnd vdd FILL
XFILL_31_NOR3X1_2 gnd vdd FILL
XFILL_33_DFFSR_117 gnd vdd FILL
XFILL_33_DFFSR_128 gnd vdd FILL
XFILL_10_NAND2X1_8 gnd vdd FILL
XFILL_2_DFFSR_141 gnd vdd FILL
XFILL_2_DFFSR_152 gnd vdd FILL
XFILL_60_DFFSR_60 gnd vdd FILL
XFILL_33_DFFSR_139 gnd vdd FILL
XFILL_2_DFFSR_163 gnd vdd FILL
XFILL_60_DFFSR_71 gnd vdd FILL
XFILL_60_DFFSR_82 gnd vdd FILL
XFILL_2_DFFSR_174 gnd vdd FILL
XFILL_60_DFFSR_93 gnd vdd FILL
XFILL_2_DFFSR_185 gnd vdd FILL
XFILL_2_DFFSR_196 gnd vdd FILL
XFILL_37_DFFSR_105 gnd vdd FILL
XFILL_37_DFFSR_116 gnd vdd FILL
XFILL_6_DFFSR_140 gnd vdd FILL
XFILL_37_DFFSR_127 gnd vdd FILL
XFILL_37_DFFSR_138 gnd vdd FILL
XFILL_26_DFFSR_4 gnd vdd FILL
XFILL_3_DFFSR_40 gnd vdd FILL
XFILL_6_DFFSR_151 gnd vdd FILL
XFILL_6_DFFSR_162 gnd vdd FILL
XFILL_3_DFFSR_51 gnd vdd FILL
XFILL_37_DFFSR_149 gnd vdd FILL
XFILL_11_NAND3X1_14 gnd vdd FILL
XFILL_10_MUX2X1_60 gnd vdd FILL
XFILL_83_DFFSR_5 gnd vdd FILL
XFILL_11_NAND3X1_25 gnd vdd FILL
XFILL_10_MUX2X1_71 gnd vdd FILL
XFILL_6_DFFSR_173 gnd vdd FILL
XFILL_3_DFFSR_62 gnd vdd FILL
XFILL_6_DFFSR_184 gnd vdd FILL
XFILL_3_DFFSR_73 gnd vdd FILL
XFILL_10_MUX2X1_82 gnd vdd FILL
XFILL_11_NAND3X1_36 gnd vdd FILL
XFILL_3_DFFSR_84 gnd vdd FILL
XFILL_11_NAND3X1_47 gnd vdd FILL
XFILL_10_MUX2X1_93 gnd vdd FILL
XFILL_6_DFFSR_195 gnd vdd FILL
XFILL_3_DFFSR_95 gnd vdd FILL
XFILL_11_NAND3X1_58 gnd vdd FILL
XFILL_2_INVX2_2 gnd vdd FILL
XFILL_11_NAND3X1_69 gnd vdd FILL
XFILL_31_CLKBUF1_14 gnd vdd FILL
XFILL_31_CLKBUF1_25 gnd vdd FILL
XFILL_31_CLKBUF1_36 gnd vdd FILL
XFILL_14_MUX2X1_70 gnd vdd FILL
XFILL_14_MUX2X1_81 gnd vdd FILL
XFILL_14_MUX2X1_92 gnd vdd FILL
XFILL_2_NOR3X1_30 gnd vdd FILL
XFILL_2_NOR3X1_41 gnd vdd FILL
XFILL_2_NOR3X1_52 gnd vdd FILL
XFILL_83_DFFSR_206 gnd vdd FILL
XFILL_34_5_1 gnd vdd FILL
XFILL_83_DFFSR_217 gnd vdd FILL
XFILL_83_DFFSR_228 gnd vdd FILL
XFILL_83_DFFSR_239 gnd vdd FILL
XFILL_33_0_0 gnd vdd FILL
XFILL_18_MUX2X1_80 gnd vdd FILL
XFILL_18_MUX2X1_91 gnd vdd FILL
XFILL_22_2 gnd vdd FILL
XFILL_6_NOR3X1_40 gnd vdd FILL
XFILL_6_NOR3X1_51 gnd vdd FILL
XFILL_48_DFFSR_8 gnd vdd FILL
XFILL_87_DFFSR_205 gnd vdd FILL
XFILL_15_1 gnd vdd FILL
XFILL_87_DFFSR_216 gnd vdd FILL
XFILL_87_DFFSR_227 gnd vdd FILL
XFILL_87_DFFSR_238 gnd vdd FILL
XFILL_22_DFFSR_160 gnd vdd FILL
XFILL_87_DFFSR_249 gnd vdd FILL
XFILL_22_DFFSR_171 gnd vdd FILL
XFILL_3_INVX1_100 gnd vdd FILL
XFILL_22_DFFSR_182 gnd vdd FILL
XFILL_3_INVX1_111 gnd vdd FILL
XFILL_3_INVX1_122 gnd vdd FILL
XFILL_22_DFFSR_193 gnd vdd FILL
XFILL_3_INVX1_133 gnd vdd FILL
XFILL_1_NAND3X1_20 gnd vdd FILL
XFILL_3_INVX1_144 gnd vdd FILL
XFILL_3_INVX1_155 gnd vdd FILL
XFILL_1_NAND3X1_31 gnd vdd FILL
XFILL_1_NAND3X1_42 gnd vdd FILL
XFILL_3_INVX1_166 gnd vdd FILL
XFILL_1_NAND3X1_53 gnd vdd FILL
XFILL_3_INVX1_177 gnd vdd FILL
XFILL_26_DFFSR_170 gnd vdd FILL
XFILL_1_NAND3X1_64 gnd vdd FILL
XFILL_5_NAND2X1_11 gnd vdd FILL
XFILL_3_INVX1_188 gnd vdd FILL
XFILL_1_NAND3X1_75 gnd vdd FILL
XFILL_5_NAND2X1_22 gnd vdd FILL
XFILL_26_DFFSR_181 gnd vdd FILL
XFILL_3_INVX1_199 gnd vdd FILL
XFILL_7_INVX1_110 gnd vdd FILL
XFILL_26_DFFSR_192 gnd vdd FILL
XFILL_5_NAND2X1_33 gnd vdd FILL
XFILL_5_NAND2X1_44 gnd vdd FILL
XFILL_1_NAND3X1_86 gnd vdd FILL
XFILL_7_INVX1_121 gnd vdd FILL
XFILL_5_NAND2X1_55 gnd vdd FILL
XFILL_1_NAND3X1_97 gnd vdd FILL
XFILL_7_INVX1_132 gnd vdd FILL
XFILL_7_INVX1_143 gnd vdd FILL
XFILL_5_NAND2X1_66 gnd vdd FILL
XFILL_7_INVX1_154 gnd vdd FILL
XFILL_5_NAND2X1_77 gnd vdd FILL
XFILL_7_INVX1_165 gnd vdd FILL
XFILL_5_NAND2X1_88 gnd vdd FILL
XINVX1_190 INVX1_190/A gnd INVX1_190/Y vdd INVX1
XFILL_7_INVX1_176 gnd vdd FILL
XFILL_7_INVX1_187 gnd vdd FILL
XFILL_7_INVX1_198 gnd vdd FILL
XFILL_13_CLKBUF1_19 gnd vdd FILL
XFILL_1_OAI22X1_6 gnd vdd FILL
XFILL_72_DFFSR_260 gnd vdd FILL
XFILL_72_DFFSR_271 gnd vdd FILL
XFILL_11_NOR2X1_104 gnd vdd FILL
XFILL_5_OAI22X1_5 gnd vdd FILL
XFILL_11_NOR2X1_115 gnd vdd FILL
XFILL_11_NOR2X1_126 gnd vdd FILL
XFILL_11_NOR2X1_137 gnd vdd FILL
XFILL_0_5_1 gnd vdd FILL
XFILL_25_5_1 gnd vdd FILL
XFILL_11_NOR2X1_148 gnd vdd FILL
XFILL_11_NOR2X1_159 gnd vdd FILL
XFILL_76_DFFSR_270 gnd vdd FILL
XFILL_24_0_0 gnd vdd FILL
XFILL_50_DFFSR_206 gnd vdd FILL
XFILL_9_AOI21X1_11 gnd vdd FILL
XFILL_9_OAI22X1_4 gnd vdd FILL
XFILL_50_DFFSR_217 gnd vdd FILL
XFILL_9_AOI21X1_22 gnd vdd FILL
XFILL_50_DFFSR_228 gnd vdd FILL
XFILL_9_AOI21X1_33 gnd vdd FILL
XFILL_50_DFFSR_239 gnd vdd FILL
XFILL_9_AOI21X1_44 gnd vdd FILL
XFILL_9_AOI21X1_55 gnd vdd FILL
XFILL_19_OAI22X1_13 gnd vdd FILL
XFILL_9_AOI21X1_66 gnd vdd FILL
XFILL_19_OAI22X1_24 gnd vdd FILL
XFILL_19_OAI22X1_35 gnd vdd FILL
XFILL_20_CLKBUF1_10 gnd vdd FILL
XFILL_9_AOI21X1_77 gnd vdd FILL
XFILL_20_CLKBUF1_21 gnd vdd FILL
XFILL_20_CLKBUF1_32 gnd vdd FILL
XFILL_54_DFFSR_205 gnd vdd FILL
XFILL_19_OAI22X1_46 gnd vdd FILL
XFILL_54_DFFSR_216 gnd vdd FILL
XFILL_54_DFFSR_227 gnd vdd FILL
XFILL_54_DFFSR_238 gnd vdd FILL
XFILL_54_DFFSR_249 gnd vdd FILL
XFILL_3_CLKBUF1_14 gnd vdd FILL
XFILL_3_CLKBUF1_25 gnd vdd FILL
XFILL_3_CLKBUF1_36 gnd vdd FILL
XFILL_81_DFFSR_105 gnd vdd FILL
XFILL_58_DFFSR_204 gnd vdd FILL
XFILL_81_DFFSR_116 gnd vdd FILL
XFILL_58_DFFSR_215 gnd vdd FILL
XFILL_81_DFFSR_127 gnd vdd FILL
XFILL_58_DFFSR_226 gnd vdd FILL
XFILL_81_DFFSR_138 gnd vdd FILL
XFILL_58_DFFSR_237 gnd vdd FILL
XFILL_81_DFFSR_149 gnd vdd FILL
XFILL_58_DFFSR_248 gnd vdd FILL
XFILL_6_BUFX2_3 gnd vdd FILL
XFILL_58_DFFSR_259 gnd vdd FILL
XFILL_85_DFFSR_104 gnd vdd FILL
XFILL_1_DFFSR_208 gnd vdd FILL
XFILL_12_OAI21X1_15 gnd vdd FILL
XFILL_1_DFFSR_219 gnd vdd FILL
XFILL_85_DFFSR_115 gnd vdd FILL
XFILL_1_NOR2X1_110 gnd vdd FILL
XFILL_85_DFFSR_126 gnd vdd FILL
XFILL_1_NOR2X1_121 gnd vdd FILL
XFILL_85_DFFSR_137 gnd vdd FILL
XFILL_12_OAI21X1_26 gnd vdd FILL
XFILL_1_NOR2X1_132 gnd vdd FILL
XFILL_8_6_1 gnd vdd FILL
XFILL_1_NOR2X1_143 gnd vdd FILL
XFILL_12_OAI21X1_37 gnd vdd FILL
XFILL_85_DFFSR_148 gnd vdd FILL
XFILL_12_OAI21X1_48 gnd vdd FILL
XFILL_7_1_0 gnd vdd FILL
XFILL_1_NOR2X1_154 gnd vdd FILL
XFILL_85_DFFSR_159 gnd vdd FILL
XFILL_1_NOR2X1_165 gnd vdd FILL
XFILL_1_NOR2X1_176 gnd vdd FILL
XFILL_1_NOR2X1_187 gnd vdd FILL
XFILL_65_DFFSR_2 gnd vdd FILL
XFILL_5_DFFSR_207 gnd vdd FILL
XFILL_8_BUFX4_11 gnd vdd FILL
XFILL_2_NAND3X1_7 gnd vdd FILL
XFILL_1_NOR2X1_198 gnd vdd FILL
XFILL_8_BUFX4_22 gnd vdd FILL
XFILL_5_DFFSR_218 gnd vdd FILL
XFILL_8_BUFX4_33 gnd vdd FILL
XFILL_5_DFFSR_229 gnd vdd FILL
XFILL_8_BUFX4_44 gnd vdd FILL
XFILL_8_BUFX4_55 gnd vdd FILL
XFILL_11_NAND2X1_80 gnd vdd FILL
XFILL_13_BUFX4_105 gnd vdd FILL
XFILL_8_BUFX4_66 gnd vdd FILL
XFILL_9_OAI22X1_30 gnd vdd FILL
XFILL_11_NAND2X1_91 gnd vdd FILL
XFILL_8_BUFX4_77 gnd vdd FILL
XFILL_9_OAI22X1_41 gnd vdd FILL
XFILL_8_BUFX4_88 gnd vdd FILL
XFILL_9_DFFSR_206 gnd vdd FILL
XFILL_8_BUFX4_99 gnd vdd FILL
XFILL_6_NAND3X1_6 gnd vdd FILL
XFILL_9_DFFSR_217 gnd vdd FILL
XFILL_9_DFFSR_228 gnd vdd FILL
XFILL_9_DFFSR_239 gnd vdd FILL
XFILL_16_5_1 gnd vdd FILL
XFILL_83_DFFSR_19 gnd vdd FILL
XFILL_15_0_0 gnd vdd FILL
XFILL_1_MUX2X1_105 gnd vdd FILL
XFILL_43_DFFSR_270 gnd vdd FILL
XNAND3X1_110 INVX1_177/A BUFX4_89/Y AND2X2_5/Y gnd NAND2X1_68/A vdd NAND3X1
XFILL_1_MUX2X1_116 gnd vdd FILL
XNAND3X1_121 DFFSR_30/Q NAND3X1_7/B NOR2X1_37/Y gnd NAND3X1_125/A vdd NAND3X1
XFILL_12_DFFSR_19 gnd vdd FILL
XNAND3X1_132 DFFSR_100/Q BUFX4_102/Y NOR2X1_37/Y gnd OAI21X1_25/C vdd NAND3X1
XFILL_1_MUX2X1_127 gnd vdd FILL
XFILL_1_MUX2X1_138 gnd vdd FILL
XFILL_1_MUX2X1_149 gnd vdd FILL
XFILL_87_DFFSR_6 gnd vdd FILL
XFILL_70_DFFSR_170 gnd vdd FILL
XFILL_2_OAI21X1_10 gnd vdd FILL
XFILL_70_DFFSR_181 gnd vdd FILL
XFILL_2_OAI21X1_21 gnd vdd FILL
XFILL_6_INVX2_3 gnd vdd FILL
XFILL_2_OAI21X1_32 gnd vdd FILL
XFILL_52_DFFSR_18 gnd vdd FILL
XFILL_70_DFFSR_192 gnd vdd FILL
XFILL_21_DFFSR_205 gnd vdd FILL
XFILL_52_DFFSR_29 gnd vdd FILL
XFILL_11_NOR2X1_18 gnd vdd FILL
XFILL_21_DFFSR_216 gnd vdd FILL
XFILL_2_OAI21X1_43 gnd vdd FILL
XFILL_11_NOR2X1_29 gnd vdd FILL
XFILL_21_DFFSR_227 gnd vdd FILL
XFILL_21_DFFSR_238 gnd vdd FILL
XFILL_21_DFFSR_249 gnd vdd FILL
XFILL_74_DFFSR_180 gnd vdd FILL
XFILL_74_DFFSR_191 gnd vdd FILL
XFILL_25_DFFSR_204 gnd vdd FILL
XFILL_25_DFFSR_215 gnd vdd FILL
XFILL_15_AOI21X1_80 gnd vdd FILL
XFILL_25_DFFSR_226 gnd vdd FILL
XFILL_4_INVX1_1 gnd vdd FILL
XFILL_25_DFFSR_237 gnd vdd FILL
XFILL_21_DFFSR_17 gnd vdd FILL
XFILL_25_DFFSR_248 gnd vdd FILL
XFILL_12_BUFX4_60 gnd vdd FILL
XFILL_21_DFFSR_28 gnd vdd FILL
XFILL_21_DFFSR_39 gnd vdd FILL
XFILL_25_DFFSR_259 gnd vdd FILL
XFILL_12_BUFX4_71 gnd vdd FILL
XFILL_78_DFFSR_190 gnd vdd FILL
XFILL_12_BUFX4_82 gnd vdd FILL
XFILL_52_DFFSR_104 gnd vdd FILL
XFILL_12_BUFX4_93 gnd vdd FILL
XFILL_29_DFFSR_203 gnd vdd FILL
XFILL_52_DFFSR_115 gnd vdd FILL
XFILL_52_DFFSR_126 gnd vdd FILL
XFILL_29_DFFSR_214 gnd vdd FILL
XFILL_29_DFFSR_225 gnd vdd FILL
XFILL_52_DFFSR_137 gnd vdd FILL
XFILL_61_DFFSR_16 gnd vdd FILL
XFILL_29_DFFSR_236 gnd vdd FILL
XFILL_52_DFFSR_148 gnd vdd FILL
XFILL_29_DFFSR_247 gnd vdd FILL
XFILL_61_DFFSR_27 gnd vdd FILL
XFILL_29_DFFSR_258 gnd vdd FILL
XFILL_52_DFFSR_159 gnd vdd FILL
XFILL_61_DFFSR_38 gnd vdd FILL
XFILL_66_4_1 gnd vdd FILL
XFILL_29_DFFSR_269 gnd vdd FILL
XFILL_61_DFFSR_49 gnd vdd FILL
XFILL_56_DFFSR_103 gnd vdd FILL
XFILL_56_DFFSR_114 gnd vdd FILL
XFILL_4_NAND3X1_19 gnd vdd FILL
XFILL_56_DFFSR_125 gnd vdd FILL
XFILL_56_DFFSR_136 gnd vdd FILL
XFILL_56_DFFSR_147 gnd vdd FILL
XFILL_56_DFFSR_158 gnd vdd FILL
XFILL_4_DFFSR_18 gnd vdd FILL
XFILL_56_DFFSR_169 gnd vdd FILL
XFILL_4_DFFSR_29 gnd vdd FILL
XFILL_30_DFFSR_15 gnd vdd FILL
XFILL_30_DFFSR_26 gnd vdd FILL
XFILL_30_DFFSR_37 gnd vdd FILL
XFILL_30_DFFSR_48 gnd vdd FILL
XFILL_6_INVX1_50 gnd vdd FILL
XFILL_30_DFFSR_59 gnd vdd FILL
XFILL_6_INVX1_61 gnd vdd FILL
XFILL_18_MUX2X1_130 gnd vdd FILL
XFILL_6_INVX1_72 gnd vdd FILL
XFILL_18_MUX2X1_141 gnd vdd FILL
XFILL_6_INVX1_83 gnd vdd FILL
XFILL_18_MUX2X1_152 gnd vdd FILL
XFILL_6_INVX1_94 gnd vdd FILL
XFILL_18_MUX2X1_163 gnd vdd FILL
XFILL_3_DFFSR_106 gnd vdd FILL
XFILL_10_DFFSR_270 gnd vdd FILL
XFILL_70_DFFSR_14 gnd vdd FILL
XFILL_3_DFFSR_117 gnd vdd FILL
XFILL_70_DFFSR_25 gnd vdd FILL
XFILL_18_MUX2X1_174 gnd vdd FILL
XFILL_18_MUX2X1_185 gnd vdd FILL
XFILL_70_DFFSR_36 gnd vdd FILL
XFILL_3_DFFSR_128 gnd vdd FILL
XFILL_70_DFFSR_47 gnd vdd FILL
XFILL_13_MUX2X1_4 gnd vdd FILL
XFILL_3_DFFSR_139 gnd vdd FILL
XFILL_70_DFFSR_58 gnd vdd FILL
XFILL_70_DFFSR_69 gnd vdd FILL
XFILL_7_DFFSR_105 gnd vdd FILL
XDFFSR_130 INVX1_165/A DFFSR_58/CLK DFFSR_91/R vdd DFFSR_130/D gnd vdd DFFSR
XFILL_7_DFFSR_116 gnd vdd FILL
XFILL_11_MUX2X1_14 gnd vdd FILL
XFILL_11_MUX2X1_25 gnd vdd FILL
XFILL_7_DFFSR_127 gnd vdd FILL
XDFFSR_141 DFFSR_141/Q CLKBUF1_8/Y DFFSR_58/R vdd DFFSR_141/D gnd vdd DFFSR
XFILL_7_DFFSR_138 gnd vdd FILL
XDFFSR_152 INVX1_150/A DFFSR_84/CLK DFFSR_82/R vdd DFFSR_152/D gnd vdd DFFSR
XFILL_11_MUX2X1_36 gnd vdd FILL
XBUFX4_4 clk gnd BUFX4_4/Y vdd BUFX4
XFILL_7_DFFSR_149 gnd vdd FILL
XFILL_4_BUFX4_70 gnd vdd FILL
XFILL_11_MUX2X1_47 gnd vdd FILL
XDFFSR_163 INVX1_148/A DFFSR_94/CLK DFFSR_99/R vdd DFFSR_163/D gnd vdd DFFSR
XFILL_2_AOI21X1_1 gnd vdd FILL
XDFFSR_174 INVX1_207/A CLKBUF1_8/Y DFFSR_89/R vdd DFFSR_174/D gnd vdd DFFSR
XFILL_11_MUX2X1_58 gnd vdd FILL
XFILL_11_MUX2X1_69 gnd vdd FILL
XFILL_4_BUFX4_81 gnd vdd FILL
XDFFSR_185 INVX1_1/A DFFSR_94/CLK DFFSR_99/R vdd DFFSR_185/D gnd vdd DFFSR
XFILL_4_BUFX4_92 gnd vdd FILL
XDFFSR_196 INVX1_137/A CLKBUF1_7/Y BUFX4_21/Y vdd DFFSR_196/D gnd vdd DFFSR
XFILL_41_DFFSR_180 gnd vdd FILL
XFILL_15_MUX2X1_13 gnd vdd FILL
XFILL_41_DFFSR_191 gnd vdd FILL
XFILL_15_MUX2X1_24 gnd vdd FILL
XFILL_15_MUX2X1_35 gnd vdd FILL
XFILL_15_MUX2X1_46 gnd vdd FILL
XFILL_15_MUX2X1_57 gnd vdd FILL
XFILL_15_MUX2X1_68 gnd vdd FILL
XFILL_15_MUX2X1_79 gnd vdd FILL
XFILL_22_MUX2X1_2 gnd vdd FILL
XFILL_3_NOR3X1_17 gnd vdd FILL
XFILL_3_NOR3X1_28 gnd vdd FILL
XFILL_45_DFFSR_190 gnd vdd FILL
XFILL_3_NOR3X1_39 gnd vdd FILL
XFILL_19_MUX2X1_12 gnd vdd FILL
XFILL_19_MUX2X1_23 gnd vdd FILL
XFILL_19_MUX2X1_34 gnd vdd FILL
XFILL_19_MUX2X1_45 gnd vdd FILL
XFILL_57_4_1 gnd vdd FILL
XFILL_6_NOR2X1_5 gnd vdd FILL
XFILL_19_MUX2X1_56 gnd vdd FILL
XFILL_19_MUX2X1_67 gnd vdd FILL
XFILL_7_NOR3X1_16 gnd vdd FILL
XFILL_19_MUX2X1_78 gnd vdd FILL
XNOR3X1_30 NOR3X1_30/A NOR3X1_30/B NOR3X1_30/C gnd NOR3X1_30/Y vdd NOR3X1
XFILL_19_MUX2X1_89 gnd vdd FILL
XFILL_7_NOR3X1_27 gnd vdd FILL
XFILL_8_MUX2X1_180 gnd vdd FILL
XNOR3X1_41 NOR3X1_41/A NOR3X1_49/B NOR3X1_6/B gnd NOR3X1_42/C vdd NOR3X1
XNOR3X1_52 NOR3X1_9/A NOR3X1_9/B NOR3X1_52/C gnd AND2X2_4/A vdd NOR3X1
XFILL_7_NOR3X1_38 gnd vdd FILL
XFILL_8_MUX2X1_191 gnd vdd FILL
XFILL_7_NOR3X1_49 gnd vdd FILL
XFILL_23_DFFSR_103 gnd vdd FILL
XFILL_23_DFFSR_114 gnd vdd FILL
XFILL_23_DFFSR_125 gnd vdd FILL
XFILL_23_DFFSR_136 gnd vdd FILL
XFILL_23_DFFSR_147 gnd vdd FILL
XFILL_23_DFFSR_158 gnd vdd FILL
XFILL_23_DFFSR_169 gnd vdd FILL
XFILL_4_INVX1_109 gnd vdd FILL
XFILL_5_MUX2X1_3 gnd vdd FILL
XFILL_27_DFFSR_102 gnd vdd FILL
XFILL_27_DFFSR_113 gnd vdd FILL
XFILL_27_DFFSR_124 gnd vdd FILL
XFILL_4_NOR2X1_109 gnd vdd FILL
XFILL_31_DFFSR_5 gnd vdd FILL
XFILL_27_DFFSR_135 gnd vdd FILL
XFILL_40_3_1 gnd vdd FILL
XFILL_10_NAND3X1_11 gnd vdd FILL
XFILL_27_DFFSR_146 gnd vdd FILL
XFILL_27_DFFSR_157 gnd vdd FILL
XFILL_10_NAND3X1_22 gnd vdd FILL
XFILL_27_DFFSR_168 gnd vdd FILL
XFILL_10_NAND3X1_33 gnd vdd FILL
XFILL_27_DFFSR_179 gnd vdd FILL
XFILL_10_NAND3X1_44 gnd vdd FILL
XFILL_69_DFFSR_3 gnd vdd FILL
XFILL_10_NAND3X1_55 gnd vdd FILL
XFILL_30_CLKBUF1_11 gnd vdd FILL
XFILL_10_NAND3X1_66 gnd vdd FILL
XFILL_30_CLKBUF1_22 gnd vdd FILL
XFILL_10_NAND3X1_77 gnd vdd FILL
XFILL_2_NOR3X1_9 gnd vdd FILL
XFILL_10_NAND3X1_88 gnd vdd FILL
XFILL_30_CLKBUF1_33 gnd vdd FILL
XFILL_10_NAND3X1_99 gnd vdd FILL
XFILL_39_DFFSR_70 gnd vdd FILL
XFILL_23_NOR3X1_14 gnd vdd FILL
XFILL_39_DFFSR_81 gnd vdd FILL
XFILL_39_DFFSR_92 gnd vdd FILL
XFILL_23_NOR3X1_25 gnd vdd FILL
XFILL_23_NOR3X1_36 gnd vdd FILL
XFILL_23_NOR3X1_47 gnd vdd FILL
XFILL_73_DFFSR_203 gnd vdd FILL
XFILL_0_DFFSR_11 gnd vdd FILL
XFILL_73_DFFSR_214 gnd vdd FILL
XFILL_0_DFFSR_22 gnd vdd FILL
XFILL_73_DFFSR_225 gnd vdd FILL
XFILL_73_DFFSR_236 gnd vdd FILL
XFILL_0_DFFSR_33 gnd vdd FILL
XFILL_73_DFFSR_247 gnd vdd FILL
XFILL_79_DFFSR_80 gnd vdd FILL
XFILL_27_NOR3X1_13 gnd vdd FILL
XFILL_73_DFFSR_258 gnd vdd FILL
XFILL_0_DFFSR_44 gnd vdd FILL
XFILL_0_DFFSR_55 gnd vdd FILL
XFILL_27_NOR3X1_24 gnd vdd FILL
XFILL_79_DFFSR_91 gnd vdd FILL
XFILL_53_DFFSR_9 gnd vdd FILL
XFILL_73_DFFSR_269 gnd vdd FILL
XFILL_0_DFFSR_66 gnd vdd FILL
XFILL_0_DFFSR_77 gnd vdd FILL
XFILL_27_NOR3X1_35 gnd vdd FILL
XFILL_77_DFFSR_202 gnd vdd FILL
XFILL_27_NOR3X1_46 gnd vdd FILL
XFILL_0_DFFSR_88 gnd vdd FILL
XFILL_77_DFFSR_213 gnd vdd FILL
XFILL_0_DFFSR_99 gnd vdd FILL
XFILL_77_DFFSR_224 gnd vdd FILL
XFILL_77_DFFSR_235 gnd vdd FILL
XFILL_1_OAI22X1_18 gnd vdd FILL
XFILL_1_OAI22X1_29 gnd vdd FILL
XFILL_77_DFFSR_246 gnd vdd FILL
XFILL_63_9 gnd vdd FILL
XFILL_77_DFFSR_257 gnd vdd FILL
XFILL_77_DFFSR_268 gnd vdd FILL
XFILL_32_CLKBUF1_9 gnd vdd FILL
XFILL_48_4_1 gnd vdd FILL
XFILL_12_DFFSR_190 gnd vdd FILL
XFILL_14_AOI22X1_11 gnd vdd FILL
XFILL_48_DFFSR_90 gnd vdd FILL
XFILL_0_NAND3X1_50 gnd vdd FILL
XFILL_0_NAND3X1_61 gnd vdd FILL
XFILL_0_NAND3X1_72 gnd vdd FILL
XFILL_0_NAND3X1_83 gnd vdd FILL
XFILL_4_NAND2X1_30 gnd vdd FILL
XFILL_4_NAND2X1_41 gnd vdd FILL
XFILL_0_NAND3X1_94 gnd vdd FILL
XFILL_4_NAND2X1_52 gnd vdd FILL
XFILL_4_NAND2X1_63 gnd vdd FILL
XFILL_4_NAND2X1_74 gnd vdd FILL
XFILL_4_NAND2X1_85 gnd vdd FILL
XFILL_4_NAND2X1_96 gnd vdd FILL
XFILL_31_3_1 gnd vdd FILL
XFILL_12_CLKBUF1_16 gnd vdd FILL
XFILL_12_CLKBUF1_27 gnd vdd FILL
XFILL_12_CLKBUF1_38 gnd vdd FILL
XFILL_10_NOR2X1_101 gnd vdd FILL
XFILL_10_NOR2X1_112 gnd vdd FILL
XFILL_10_NOR2X1_123 gnd vdd FILL
XFILL_10_NOR2X1_134 gnd vdd FILL
XFILL_10_NOR2X1_145 gnd vdd FILL
XFILL_10_NOR2X1_156 gnd vdd FILL
XFILL_10_NOR2X1_167 gnd vdd FILL
XFILL_10_NOR2X1_178 gnd vdd FILL
XFILL_40_DFFSR_203 gnd vdd FILL
XFILL_10_NOR2X1_189 gnd vdd FILL
XFILL_40_DFFSR_214 gnd vdd FILL
XFILL_2_OAI21X1_4 gnd vdd FILL
XFILL_40_DFFSR_225 gnd vdd FILL
XFILL_8_AOI21X1_30 gnd vdd FILL
XFILL_40_DFFSR_236 gnd vdd FILL
XFILL_8_AOI21X1_41 gnd vdd FILL
XFILL_40_DFFSR_247 gnd vdd FILL
XFILL_8_AOI21X1_52 gnd vdd FILL
XFILL_40_DFFSR_258 gnd vdd FILL
XFILL_18_OAI22X1_10 gnd vdd FILL
XFILL_8_AOI21X1_63 gnd vdd FILL
XFILL_40_DFFSR_269 gnd vdd FILL
XNAND3X1_7 DFFSR_31/Q NAND3X1_7/B NOR2X1_37/Y gnd NAND3X1_8/A vdd NAND3X1
XFILL_18_OAI22X1_21 gnd vdd FILL
XFILL_8_AOI21X1_74 gnd vdd FILL
XFILL_18_OAI22X1_32 gnd vdd FILL
XFILL_44_DFFSR_202 gnd vdd FILL
XFILL_18_OAI22X1_43 gnd vdd FILL
XFILL_6_OAI21X1_3 gnd vdd FILL
XFILL_44_DFFSR_213 gnd vdd FILL
XFILL_39_4_1 gnd vdd FILL
XFILL_44_DFFSR_224 gnd vdd FILL
XFILL_44_DFFSR_235 gnd vdd FILL
XFILL_3_NOR2X1_50 gnd vdd FILL
XFILL_44_DFFSR_246 gnd vdd FILL
XFILL_2_CLKBUF1_11 gnd vdd FILL
XFILL_3_NOR2X1_61 gnd vdd FILL
XFILL_44_DFFSR_257 gnd vdd FILL
XFILL_13_BUFX4_16 gnd vdd FILL
XFILL_3_NOR2X1_72 gnd vdd FILL
XFILL_2_CLKBUF1_22 gnd vdd FILL
XFILL_44_DFFSR_268 gnd vdd FILL
XFILL_13_BUFX4_27 gnd vdd FILL
XFILL_3_NOR2X1_83 gnd vdd FILL
XFILL_3_NOR2X1_94 gnd vdd FILL
XFILL_2_CLKBUF1_33 gnd vdd FILL
XFILL_13_BUFX4_38 gnd vdd FILL
XFILL_48_DFFSR_201 gnd vdd FILL
XFILL_71_DFFSR_102 gnd vdd FILL
XFILL_48_DFFSR_212 gnd vdd FILL
XFILL_13_BUFX4_49 gnd vdd FILL
XFILL_71_DFFSR_113 gnd vdd FILL
XFILL_10_MUX2X1_107 gnd vdd FILL
XFILL_71_DFFSR_124 gnd vdd FILL
XFILL_10_MUX2X1_118 gnd vdd FILL
XFILL_10_MUX2X1_129 gnd vdd FILL
XFILL_71_DFFSR_135 gnd vdd FILL
XFILL_48_DFFSR_223 gnd vdd FILL
XFILL_48_DFFSR_234 gnd vdd FILL
XFILL_71_DFFSR_146 gnd vdd FILL
XFILL_7_NOR2X1_60 gnd vdd FILL
XFILL_48_DFFSR_245 gnd vdd FILL
XFILL_71_DFFSR_157 gnd vdd FILL
XFILL_48_DFFSR_256 gnd vdd FILL
XFILL_48_DFFSR_267 gnd vdd FILL
XFILL_7_NOR2X1_71 gnd vdd FILL
XFILL_71_DFFSR_168 gnd vdd FILL
XFILL_71_DFFSR_179 gnd vdd FILL
XFILL_7_NOR2X1_82 gnd vdd FILL
XFILL_7_NOR2X1_93 gnd vdd FILL
XFILL_75_DFFSR_101 gnd vdd FILL
XFILL_11_OAI21X1_12 gnd vdd FILL
XFILL_75_DFFSR_112 gnd vdd FILL
XFILL_75_DFFSR_123 gnd vdd FILL
XFILL_75_DFFSR_134 gnd vdd FILL
XFILL_11_OAI21X1_23 gnd vdd FILL
XFILL_22_3_1 gnd vdd FILL
XFILL_0_DFFSR_4 gnd vdd FILL
XFILL_75_DFFSR_145 gnd vdd FILL
XFILL_0_NOR2X1_140 gnd vdd FILL
XFILL_11_OAI21X1_34 gnd vdd FILL
XFILL_11_OAI21X1_45 gnd vdd FILL
XFILL_75_DFFSR_156 gnd vdd FILL
XFILL_0_NOR2X1_151 gnd vdd FILL
XFILL_13_DFFSR_2 gnd vdd FILL
XFILL_0_NOR2X1_162 gnd vdd FILL
XFILL_75_DFFSR_167 gnd vdd FILL
XFILL_70_DFFSR_3 gnd vdd FILL
XFILL_75_DFFSR_178 gnd vdd FILL
XFILL_0_NOR2X1_173 gnd vdd FILL
XFILL_79_DFFSR_100 gnd vdd FILL
XFILL_0_NOR2X1_184 gnd vdd FILL
XFILL_75_DFFSR_189 gnd vdd FILL
XFILL_0_NOR2X1_195 gnd vdd FILL
XFILL_79_DFFSR_111 gnd vdd FILL
XFILL_79_DFFSR_122 gnd vdd FILL
XFILL_79_DFFSR_133 gnd vdd FILL
XFILL_79_DFFSR_144 gnd vdd FILL
XFILL_79_DFFSR_155 gnd vdd FILL
XFILL_7_INVX1_17 gnd vdd FILL
XFILL_7_INVX1_28 gnd vdd FILL
XFILL_79_DFFSR_166 gnd vdd FILL
XFILL_79_DFFSR_177 gnd vdd FILL
XFILL_7_INVX1_39 gnd vdd FILL
XFILL_79_DFFSR_188 gnd vdd FILL
XFILL_79_DFFSR_199 gnd vdd FILL
XBUFX2_1 BUFX2_1/A gnd dout[1] vdd BUFX2
XFILL_0_MUX2X1_102 gnd vdd FILL
XFILL_0_MUX2X1_113 gnd vdd FILL
XFILL_3_NAND2X1_5 gnd vdd FILL
XFILL_0_MUX2X1_124 gnd vdd FILL
XFILL_0_MUX2X1_135 gnd vdd FILL
XFILL_0_MUX2X1_146 gnd vdd FILL
XFILL_35_DFFSR_6 gnd vdd FILL
XFILL_5_BUFX4_15 gnd vdd FILL
XFILL_0_MUX2X1_157 gnd vdd FILL
XFILL_5_BUFX4_26 gnd vdd FILL
XFILL_0_MUX2X1_168 gnd vdd FILL
XFILL_5_BUFX4_37 gnd vdd FILL
XFILL_5_BUFX4_48 gnd vdd FILL
XFILL_0_MUX2X1_179 gnd vdd FILL
XFILL_5_BUFX4_59 gnd vdd FILL
XFILL_5_4_1 gnd vdd FILL
XFILL_7_NAND2X1_4 gnd vdd FILL
XFILL_11_DFFSR_202 gnd vdd FILL
XFILL_1_OAI21X1_40 gnd vdd FILL
XFILL_11_DFFSR_213 gnd vdd FILL
XFILL_11_DFFSR_224 gnd vdd FILL
XFILL_11_DFFSR_235 gnd vdd FILL
XFILL_11_DFFSR_246 gnd vdd FILL
XFILL_3_MUX2X1_90 gnd vdd FILL
XFILL_11_DFFSR_257 gnd vdd FILL
XFILL_11_DFFSR_268 gnd vdd FILL
XFILL_15_DFFSR_201 gnd vdd FILL
XFILL_15_DFFSR_212 gnd vdd FILL
XFILL_12_NAND3X1_1 gnd vdd FILL
XFILL_15_DFFSR_223 gnd vdd FILL
XFILL_15_DFFSR_234 gnd vdd FILL
XFILL_15_DFFSR_245 gnd vdd FILL
XFILL_15_DFFSR_256 gnd vdd FILL
XFILL_15_DFFSR_267 gnd vdd FILL
XFILL_13_3_1 gnd vdd FILL
XFILL_42_DFFSR_101 gnd vdd FILL
XFILL_19_DFFSR_200 gnd vdd FILL
XFILL_12_AND2X2_3 gnd vdd FILL
XFILL_19_DFFSR_211 gnd vdd FILL
XFILL_42_DFFSR_112 gnd vdd FILL
XFILL_42_DFFSR_123 gnd vdd FILL
XFILL_42_DFFSR_134 gnd vdd FILL
XFILL_19_DFFSR_222 gnd vdd FILL
XINVX2_1 INVX2_1/A gnd OR2X2_1/A vdd INVX2
XFILL_19_DFFSR_233 gnd vdd FILL
XFILL_42_DFFSR_145 gnd vdd FILL
XFILL_19_DFFSR_244 gnd vdd FILL
XFILL_42_DFFSR_156 gnd vdd FILL
XFILL_19_DFFSR_255 gnd vdd FILL
XFILL_42_DFFSR_167 gnd vdd FILL
XFILL_19_DFFSR_266 gnd vdd FILL
XFILL_42_DFFSR_178 gnd vdd FILL
XFILL_42_DFFSR_189 gnd vdd FILL
XFILL_46_DFFSR_100 gnd vdd FILL
XFILL_46_DFFSR_111 gnd vdd FILL
XAOI21X1_1 BUFX4_72/Y AOI21X1_1/B AOI21X1_1/C gnd DFFSR_181/D vdd AOI21X1
XFILL_3_NAND3X1_16 gnd vdd FILL
XFILL_46_DFFSR_122 gnd vdd FILL
XFILL_7_AOI21X1_9 gnd vdd FILL
XFILL_46_DFFSR_133 gnd vdd FILL
XFILL_3_NAND3X1_27 gnd vdd FILL
XFILL_46_DFFSR_144 gnd vdd FILL
XFILL_3_NAND3X1_38 gnd vdd FILL
XFILL_46_DFFSR_155 gnd vdd FILL
XFILL_3_NAND3X1_49 gnd vdd FILL
XFILL_46_DFFSR_166 gnd vdd FILL
XFILL_46_DFFSR_177 gnd vdd FILL
XFILL_7_NAND2X1_18 gnd vdd FILL
XFILL_46_DFFSR_188 gnd vdd FILL
XFILL_7_NAND2X1_29 gnd vdd FILL
XFILL_46_DFFSR_199 gnd vdd FILL
XMUX2X1_170 BUFX4_80/Y INVX1_215/Y NOR2X1_165/Y gnd DFFSR_67/D vdd MUX2X1
XFILL_12_AOI22X1_6 gnd vdd FILL
XMUX2X1_181 BUFX4_74/Y INVX1_226/Y NOR2X1_167/Y gnd DFFSR_61/D vdd MUX2X1
XMUX2X1_192 MUX2X1_8/A NOR3X1_5/A MUX2X1_3/S gnd DFFSR_45/D vdd MUX2X1
XFILL_5_4 gnd vdd FILL
XFILL_17_MUX2X1_160 gnd vdd FILL
XFILL_17_MUX2X1_171 gnd vdd FILL
XFILL_17_MUX2X1_182 gnd vdd FILL
XFILL_17_MUX2X1_193 gnd vdd FILL
XFILL_16_AOI22X1_5 gnd vdd FILL
XFILL_54_5 gnd vdd FILL
XFILL_64_7_2 gnd vdd FILL
XFILL_3_INVX1_10 gnd vdd FILL
XFILL_3_INVX1_21 gnd vdd FILL
XFILL_63_2_1 gnd vdd FILL
XFILL_3_INVX1_32 gnd vdd FILL
XFILL_3_INVX1_43 gnd vdd FILL
XFILL_4_AND2X2_2 gnd vdd FILL
XFILL_3_INVX1_54 gnd vdd FILL
XFILL_3_INVX1_65 gnd vdd FILL
XFILL_3_INVX1_76 gnd vdd FILL
XFILL_49_DFFSR_13 gnd vdd FILL
XFILL_3_INVX1_87 gnd vdd FILL
XFILL_49_DFFSR_24 gnd vdd FILL
XFILL_49_DFFSR_35 gnd vdd FILL
XFILL_3_INVX1_98 gnd vdd FILL
XFILL_49_DFFSR_46 gnd vdd FILL
XFILL_49_DFFSR_57 gnd vdd FILL
XFILL_49_DFFSR_68 gnd vdd FILL
XFILL_10_MUX2X1_8 gnd vdd FILL
XFILL_49_DFFSR_79 gnd vdd FILL
XFILL_22_CLKBUF1_17 gnd vdd FILL
XFILL_22_CLKBUF1_28 gnd vdd FILL
XFILL_1_BUFX4_30 gnd vdd FILL
XFILL_22_CLKBUF1_39 gnd vdd FILL
XFILL_1_BUFX4_41 gnd vdd FILL
XFILL_18_DFFSR_12 gnd vdd FILL
XFILL_1_BUFX4_52 gnd vdd FILL
XFILL_1_BUFX4_63 gnd vdd FILL
XFILL_18_DFFSR_23 gnd vdd FILL
XFILL_18_DFFSR_34 gnd vdd FILL
XFILL_1_BUFX4_74 gnd vdd FILL
XFILL_18_DFFSR_45 gnd vdd FILL
XFILL_18_DFFSR_56 gnd vdd FILL
XFILL_1_BUFX4_85 gnd vdd FILL
XFILL_1_BUFX4_96 gnd vdd FILL
XFILL_18_DFFSR_67 gnd vdd FILL
XFILL_13_DFFSR_100 gnd vdd FILL
XFILL_13_DFFSR_111 gnd vdd FILL
XFILL_18_DFFSR_78 gnd vdd FILL
XFILL_13_DFFSR_122 gnd vdd FILL
XFILL_18_DFFSR_89 gnd vdd FILL
XFILL_0_AOI21X1_18 gnd vdd FILL
XFILL_13_DFFSR_133 gnd vdd FILL
XFILL_13_DFFSR_144 gnd vdd FILL
XFILL_58_DFFSR_11 gnd vdd FILL
XFILL_0_AOI21X1_29 gnd vdd FILL
XFILL_58_DFFSR_22 gnd vdd FILL
XFILL_13_DFFSR_155 gnd vdd FILL
XFILL_13_DFFSR_166 gnd vdd FILL
XFILL_58_DFFSR_33 gnd vdd FILL
XFILL_29_NOR3X1_8 gnd vdd FILL
XFILL_2_CLKBUF1_9 gnd vdd FILL
XFILL_13_DFFSR_177 gnd vdd FILL
XFILL_58_DFFSR_44 gnd vdd FILL
XFILL_58_DFFSR_55 gnd vdd FILL
XFILL_13_DFFSR_188 gnd vdd FILL
XFILL_58_DFFSR_66 gnd vdd FILL
XFILL_58_DFFSR_77 gnd vdd FILL
XFILL_17_DFFSR_110 gnd vdd FILL
XFILL_13_DFFSR_199 gnd vdd FILL
XFILL_3_NOR2X1_106 gnd vdd FILL
XFILL_17_DFFSR_121 gnd vdd FILL
XFILL_17_DFFSR_132 gnd vdd FILL
XFILL_58_DFFSR_88 gnd vdd FILL
XFILL_3_NOR2X1_117 gnd vdd FILL
XFILL_4_DFFSR_5 gnd vdd FILL
XFILL_17_DFFSR_143 gnd vdd FILL
XFILL_58_DFFSR_99 gnd vdd FILL
XFILL_3_NOR2X1_128 gnd vdd FILL
XFILL_3_NOR2X1_139 gnd vdd FILL
XFILL_17_DFFSR_3 gnd vdd FILL
XFILL_17_DFFSR_154 gnd vdd FILL
XFILL_17_DFFSR_165 gnd vdd FILL
XFILL_74_DFFSR_4 gnd vdd FILL
XFILL_3_NOR2X1_9 gnd vdd FILL
XFILL_6_CLKBUF1_8 gnd vdd FILL
XFILL_17_DFFSR_176 gnd vdd FILL
XFILL_17_DFFSR_187 gnd vdd FILL
XFILL_27_DFFSR_10 gnd vdd FILL
XFILL_27_DFFSR_21 gnd vdd FILL
XFILL_17_DFFSR_198 gnd vdd FILL
XFILL_27_DFFSR_32 gnd vdd FILL
XFILL_27_DFFSR_43 gnd vdd FILL
XFILL_27_DFFSR_54 gnd vdd FILL
XFILL_27_DFFSR_65 gnd vdd FILL
XFILL_27_DFFSR_76 gnd vdd FILL
XFILL_2_BUFX4_103 gnd vdd FILL
XFILL_55_7_2 gnd vdd FILL
XFILL_27_DFFSR_87 gnd vdd FILL
XFILL_13_NOR3X1_11 gnd vdd FILL
XFILL_27_DFFSR_98 gnd vdd FILL
XFILL_13_NOR3X1_22 gnd vdd FILL
XFILL_54_2_1 gnd vdd FILL
XFILL_67_DFFSR_20 gnd vdd FILL
XFILL_13_NOR3X1_33 gnd vdd FILL
XFILL_67_DFFSR_31 gnd vdd FILL
XFILL_63_DFFSR_200 gnd vdd FILL
XFILL_13_NOR3X1_44 gnd vdd FILL
XFILL_67_DFFSR_42 gnd vdd FILL
XFILL_63_DFFSR_211 gnd vdd FILL
XFILL_20_MUX2X1_108 gnd vdd FILL
XFILL_2_MUX2X1_7 gnd vdd FILL
XFILL_20_MUX2X1_119 gnd vdd FILL
XFILL_67_DFFSR_53 gnd vdd FILL
XFILL_63_DFFSR_222 gnd vdd FILL
XFILL_6_BUFX4_102 gnd vdd FILL
XFILL_67_DFFSR_64 gnd vdd FILL
XFILL_63_DFFSR_233 gnd vdd FILL
XFILL_67_DFFSR_75 gnd vdd FILL
XFILL_67_DFFSR_86 gnd vdd FILL
XFILL_63_DFFSR_244 gnd vdd FILL
XFILL_17_NOR3X1_10 gnd vdd FILL
XFILL_63_DFFSR_255 gnd vdd FILL
XFILL_67_DFFSR_97 gnd vdd FILL
XFILL_17_NOR3X1_21 gnd vdd FILL
XFILL_63_DFFSR_266 gnd vdd FILL
XFILL_17_NOR3X1_32 gnd vdd FILL
XFILL_17_NOR3X1_43 gnd vdd FILL
XFILL_67_DFFSR_210 gnd vdd FILL
XFILL_39_DFFSR_7 gnd vdd FILL
XFILL_8_NOR2X1_206 gnd vdd FILL
XFILL_67_DFFSR_221 gnd vdd FILL
XFILL_0_OAI22X1_15 gnd vdd FILL
XFILL_36_DFFSR_30 gnd vdd FILL
XFILL_67_DFFSR_232 gnd vdd FILL
XFILL_67_DFFSR_243 gnd vdd FILL
XFILL_36_DFFSR_41 gnd vdd FILL
XFILL_0_OAI22X1_26 gnd vdd FILL
XFILL_67_DFFSR_254 gnd vdd FILL
XFILL_0_OAI22X1_37 gnd vdd FILL
XFILL_36_DFFSR_52 gnd vdd FILL
XFILL_67_DFFSR_265 gnd vdd FILL
XFILL_0_OAI22X1_48 gnd vdd FILL
XFILL_36_DFFSR_63 gnd vdd FILL
XFILL_22_CLKBUF1_6 gnd vdd FILL
XFILL_4_OAI21X1_17 gnd vdd FILL
XFILL_36_DFFSR_74 gnd vdd FILL
XFILL_4_OAI21X1_28 gnd vdd FILL
XFILL_36_DFFSR_85 gnd vdd FILL
XAOI21X1_20 MUX2X1_2/A NOR2X1_161/B NOR2X1_161/Y gnd DFFSR_84/D vdd AOI21X1
XFILL_36_DFFSR_96 gnd vdd FILL
XFILL_4_OAI21X1_39 gnd vdd FILL
XFILL_0_NOR2X1_16 gnd vdd FILL
XFILL_0_NOR2X1_27 gnd vdd FILL
XAOI21X1_31 BUFX4_65/Y NOR2X1_190/B NOR2X1_188/Y gnd DFFSR_20/D vdd AOI21X1
XAOI21X1_42 BUFX4_97/Y NOR2X1_202/B NOR2X1_202/Y gnd DFFSR_9/D vdd AOI21X1
XFILL_0_NOR2X1_38 gnd vdd FILL
XAOI21X1_53 BUFX4_97/Y NOR2X1_12/B NOR2X1_12/Y gnd DFFSR_266/D vdd AOI21X1
XFILL_76_DFFSR_40 gnd vdd FILL
XFILL_0_NOR2X1_49 gnd vdd FILL
XFILL_76_DFFSR_51 gnd vdd FILL
XAOI21X1_64 OAI21X1_42/Y NAND3X1_43/B DFFSR_1/D gnd AND2X2_6/B vdd AOI21X1
XFILL_76_DFFSR_62 gnd vdd FILL
XAOI21X1_75 NAND3X1_31/Y BUFX2_9/A AOI22X1_3/A gnd AOI22X1_2/D vdd AOI21X1
XFILL_26_CLKBUF1_5 gnd vdd FILL
XFILL_76_DFFSR_73 gnd vdd FILL
XFILL_76_DFFSR_84 gnd vdd FILL
XOAI21X1_4 OAI21X1_4/A OAI21X1_4/B OAI21X1_4/C gnd OAI21X1_4/Y vdd OAI21X1
XFILL_76_DFFSR_95 gnd vdd FILL
XFILL_3_NAND2X1_60 gnd vdd FILL
XFILL_4_NOR2X1_15 gnd vdd FILL
XFILL_4_NOR2X1_26 gnd vdd FILL
XFILL_3_NAND2X1_71 gnd vdd FILL
XFILL_11_BUFX4_3 gnd vdd FILL
XFILL_4_NOR2X1_37 gnd vdd FILL
XFILL_3_NAND2X1_82 gnd vdd FILL
XFILL_4_NOR2X1_48 gnd vdd FILL
XFILL_3_NAND2X1_93 gnd vdd FILL
XFILL_4_NOR2X1_59 gnd vdd FILL
XFILL_16_NOR3X1_3 gnd vdd FILL
XFILL_11_CLKBUF1_13 gnd vdd FILL
XFILL_11_CLKBUF1_24 gnd vdd FILL
XFILL_8_NOR2X1_14 gnd vdd FILL
XFILL_45_DFFSR_50 gnd vdd FILL
XFILL_8_NOR2X1_25 gnd vdd FILL
XFILL_11_CLKBUF1_35 gnd vdd FILL
XFILL_45_DFFSR_61 gnd vdd FILL
XFILL_8_NOR2X1_36 gnd vdd FILL
XFILL_45_DFFSR_72 gnd vdd FILL
XFILL_8_NOR2X1_47 gnd vdd FILL
XFILL_45_DFFSR_83 gnd vdd FILL
XFILL_8_NOR2X1_58 gnd vdd FILL
XFILL_45_DFFSR_94 gnd vdd FILL
XFILL_12_OAI22X1_9 gnd vdd FILL
XFILL_8_NOR2X1_69 gnd vdd FILL
XFILL_46_7_2 gnd vdd FILL
XFILL_85_DFFSR_60 gnd vdd FILL
XFILL_85_DFFSR_71 gnd vdd FILL
XFILL_85_DFFSR_82 gnd vdd FILL
XFILL_45_2_1 gnd vdd FILL
XFILL_16_OAI22X1_8 gnd vdd FILL
XFILL_85_DFFSR_93 gnd vdd FILL
XFILL_14_DFFSR_60 gnd vdd FILL
XFILL_14_DFFSR_71 gnd vdd FILL
XFILL_14_DFFSR_82 gnd vdd FILL
XFILL_14_DFFSR_93 gnd vdd FILL
XFILL_30_DFFSR_200 gnd vdd FILL
XFILL_30_DFFSR_211 gnd vdd FILL
XFILL_30_DFFSR_222 gnd vdd FILL
XFILL_25_NOR3X1_1 gnd vdd FILL
XFILL_26_9 gnd vdd FILL
XFILL_30_DFFSR_233 gnd vdd FILL
XFILL_30_DFFSR_244 gnd vdd FILL
XFILL_30_DFFSR_255 gnd vdd FILL
XOAI22X1_50 INVX1_183/Y OAI22X1_50/B INVX1_179/Y OAI22X1_50/D gnd NOR2X1_49/B vdd
+ OAI22X1
XFILL_7_AOI21X1_60 gnd vdd FILL
XFILL_54_DFFSR_70 gnd vdd FILL
XFILL_7_AOI21X1_71 gnd vdd FILL
XFILL_54_DFFSR_81 gnd vdd FILL
XFILL_30_DFFSR_266 gnd vdd FILL
XFILL_54_DFFSR_92 gnd vdd FILL
XFILL_17_OAI22X1_40 gnd vdd FILL
XFILL_17_OAI22X1_51 gnd vdd FILL
XFILL_34_DFFSR_210 gnd vdd FILL
XFILL_34_DFFSR_221 gnd vdd FILL
XFILL_34_DFFSR_232 gnd vdd FILL
XFILL_34_DFFSR_243 gnd vdd FILL
XFILL_34_DFFSR_254 gnd vdd FILL
XFILL_34_DFFSR_265 gnd vdd FILL
XFILL_0_MUX2X1_12 gnd vdd FILL
XFILL_1_CLKBUF1_30 gnd vdd FILL
XFILL_0_MUX2X1_23 gnd vdd FILL
XFILL_1_CLKBUF1_41 gnd vdd FILL
XFILL_0_MUX2X1_34 gnd vdd FILL
XFILL_1_INVX8_3 gnd vdd FILL
XFILL_0_MUX2X1_45 gnd vdd FILL
XFILL_61_DFFSR_110 gnd vdd FILL
XFILL_38_DFFSR_220 gnd vdd FILL
XFILL_61_DFFSR_121 gnd vdd FILL
XFILL_23_DFFSR_80 gnd vdd FILL
XFILL_14_INVX8_1 gnd vdd FILL
XFILL_61_DFFSR_132 gnd vdd FILL
XFILL_0_MUX2X1_56 gnd vdd FILL
XFILL_61_DFFSR_143 gnd vdd FILL
XFILL_23_DFFSR_91 gnd vdd FILL
XFILL_38_DFFSR_231 gnd vdd FILL
XFILL_0_MUX2X1_67 gnd vdd FILL
XFILL_0_MUX2X1_78 gnd vdd FILL
XFILL_38_DFFSR_242 gnd vdd FILL
XFILL_8_NOR3X1_2 gnd vdd FILL
XFILL_61_DFFSR_154 gnd vdd FILL
XFILL_38_DFFSR_253 gnd vdd FILL
XFILL_0_MUX2X1_89 gnd vdd FILL
XFILL_61_DFFSR_165 gnd vdd FILL
XFILL_38_DFFSR_264 gnd vdd FILL
XFILL_38_DFFSR_275 gnd vdd FILL
XFILL_4_MUX2X1_11 gnd vdd FILL
XFILL_61_DFFSR_176 gnd vdd FILL
XFILL_4_MUX2X1_22 gnd vdd FILL
XFILL_61_DFFSR_187 gnd vdd FILL
XFILL_4_MUX2X1_33 gnd vdd FILL
XFILL_61_DFFSR_198 gnd vdd FILL
XFILL_4_MUX2X1_44 gnd vdd FILL
XFILL_10_OAI21X1_20 gnd vdd FILL
XFILL_65_DFFSR_120 gnd vdd FILL
XFILL_4_MUX2X1_55 gnd vdd FILL
XFILL_65_DFFSR_131 gnd vdd FILL
XFILL_63_DFFSR_90 gnd vdd FILL
XFILL_65_DFFSR_142 gnd vdd FILL
XFILL_4_MUX2X1_66 gnd vdd FILL
XFILL_10_OAI21X1_31 gnd vdd FILL
XFILL_4_MUX2X1_77 gnd vdd FILL
XFILL_65_DFFSR_153 gnd vdd FILL
XFILL_3_1 gnd vdd FILL
XFILL_10_OAI21X1_42 gnd vdd FILL
XFILL_4_MUX2X1_88 gnd vdd FILL
XFILL_4_MUX2X1_99 gnd vdd FILL
XFILL_8_MUX2X1_10 gnd vdd FILL
XFILL_65_DFFSR_164 gnd vdd FILL
XFILL_65_DFFSR_175 gnd vdd FILL
XFILL_8_MUX2X1_21 gnd vdd FILL
XFILL_65_DFFSR_186 gnd vdd FILL
XFILL_65_DFFSR_197 gnd vdd FILL
XFILL_8_MUX2X1_32 gnd vdd FILL
XFILL_56_DFFSR_1 gnd vdd FILL
XFILL_8_MUX2X1_43 gnd vdd FILL
XFILL_8_MUX2X1_54 gnd vdd FILL
XFILL_69_DFFSR_130 gnd vdd FILL
XFILL_6_DFFSR_70 gnd vdd FILL
XFILL_8_MUX2X1_65 gnd vdd FILL
XFILL_69_DFFSR_141 gnd vdd FILL
XFILL_69_DFFSR_152 gnd vdd FILL
XFILL_8_MUX2X1_76 gnd vdd FILL
XFILL_6_DFFSR_81 gnd vdd FILL
XFILL_8_MUX2X1_87 gnd vdd FILL
XFILL_6_DFFSR_92 gnd vdd FILL
XFILL_37_7_2 gnd vdd FILL
XFILL_69_DFFSR_163 gnd vdd FILL
XFILL_8_MUX2X1_98 gnd vdd FILL
XFILL_69_DFFSR_174 gnd vdd FILL
XFILL_69_DFFSR_185 gnd vdd FILL
XFILL_45_1 gnd vdd FILL
XFILL_36_2_1 gnd vdd FILL
XFILL_69_DFFSR_196 gnd vdd FILL
XFILL_47_DFFSR_109 gnd vdd FILL
XFILL_20_MUX2X1_20 gnd vdd FILL
XFILL_20_MUX2X1_31 gnd vdd FILL
XFILL_40_DFFSR_7 gnd vdd FILL
XFILL_8_DFFSR_6 gnd vdd FILL
XFILL_20_MUX2X1_42 gnd vdd FILL
XFILL_20_MUX2X1_53 gnd vdd FILL
XFILL_12_NAND3X1_18 gnd vdd FILL
XFILL_20_MUX2X1_64 gnd vdd FILL
XFILL_20_MUX2X1_75 gnd vdd FILL
XFILL_12_NAND3X1_29 gnd vdd FILL
XFILL_20_6_2 gnd vdd FILL
XFILL_78_DFFSR_5 gnd vdd FILL
XFILL_20_MUX2X1_86 gnd vdd FILL
XFILL_20_MUX2X1_97 gnd vdd FILL
XFILL_32_CLKBUF1_18 gnd vdd FILL
XFILL_32_CLKBUF1_29 gnd vdd FILL
XFILL_2_BUFX4_19 gnd vdd FILL
XFILL_32_DFFSR_120 gnd vdd FILL
XFILL_32_DFFSR_131 gnd vdd FILL
XFILL_32_DFFSR_142 gnd vdd FILL
XFILL_32_DFFSR_153 gnd vdd FILL
XFILL_32_DFFSR_164 gnd vdd FILL
XFILL_32_DFFSR_175 gnd vdd FILL
XFILL_32_DFFSR_186 gnd vdd FILL
XFILL_32_DFFSR_197 gnd vdd FILL
XFILL_2_NAND3X1_13 gnd vdd FILL
XFILL_28_7_2 gnd vdd FILL
XFILL_36_DFFSR_130 gnd vdd FILL
XFILL_3_7_2 gnd vdd FILL
XFILL_2_NAND3X1_24 gnd vdd FILL
XFILL_2_NAND3X1_35 gnd vdd FILL
XFILL_36_DFFSR_141 gnd vdd FILL
XFILL_36_DFFSR_152 gnd vdd FILL
XFILL_27_2_1 gnd vdd FILL
XFILL_2_2_1 gnd vdd FILL
XFILL_2_NAND3X1_46 gnd vdd FILL
XFILL_2_NAND3X1_57 gnd vdd FILL
XFILL_36_DFFSR_163 gnd vdd FILL
XFILL_6_NAND2X1_15 gnd vdd FILL
XFILL_36_DFFSR_174 gnd vdd FILL
XFILL_2_NAND3X1_68 gnd vdd FILL
XFILL_6_NAND2X1_26 gnd vdd FILL
XFILL_2_NAND3X1_79 gnd vdd FILL
XFILL_36_DFFSR_185 gnd vdd FILL
XFILL_6_NAND2X1_37 gnd vdd FILL
XFILL_36_DFFSR_196 gnd vdd FILL
XFILL_6_NAND2X1_48 gnd vdd FILL
XFILL_2_BUFX4_6 gnd vdd FILL
XFILL_6_NAND2X1_59 gnd vdd FILL
XFILL_15_BUFX4_4 gnd vdd FILL
XMUX2X1_8 MUX2X1_8/A NOR3X1_6/A MUX2X1_9/S gnd MUX2X1_8/Y vdd MUX2X1
XFILL_14_DFFSR_109 gnd vdd FILL
XFILL_16_MUX2X1_190 gnd vdd FILL
XFILL_11_6_2 gnd vdd FILL
XFILL_82_DFFSR_220 gnd vdd FILL
XFILL_10_1_1 gnd vdd FILL
XFILL_82_DFFSR_231 gnd vdd FILL
XFILL_82_DFFSR_242 gnd vdd FILL
XFILL_82_DFFSR_253 gnd vdd FILL
XFILL_82_DFFSR_264 gnd vdd FILL
XFILL_82_DFFSR_275 gnd vdd FILL
XFILL_18_DFFSR_108 gnd vdd FILL
XFILL_18_DFFSR_119 gnd vdd FILL
XFILL_13_AOI21X1_4 gnd vdd FILL
XFILL_86_DFFSR_230 gnd vdd FILL
XCLKBUF1_9 BUFX4_95/Y gnd DFFSR_6/CLK vdd CLKBUF1
XFILL_86_DFFSR_241 gnd vdd FILL
XFILL_86_DFFSR_252 gnd vdd FILL
XFILL_86_DFFSR_263 gnd vdd FILL
XFILL_86_DFFSR_274 gnd vdd FILL
XFILL_37_DFFSR_19 gnd vdd FILL
XFILL_2_INVX1_180 gnd vdd FILL
XFILL_2_INVX1_191 gnd vdd FILL
XFILL_77_DFFSR_18 gnd vdd FILL
XFILL_77_DFFSR_29 gnd vdd FILL
XFILL_21_CLKBUF1_14 gnd vdd FILL
XFILL_21_CLKBUF1_25 gnd vdd FILL
XFILL_64_DFFSR_209 gnd vdd FILL
XFILL_21_CLKBUF1_36 gnd vdd FILL
XBUFX4_103 BUFX4_2/A gnd BUFX4_103/Y vdd BUFX4
XFILL_0_INVX1_14 gnd vdd FILL
XFILL_0_INVX1_25 gnd vdd FILL
XFILL_0_INVX1_36 gnd vdd FILL
XFILL_6_INVX1_190 gnd vdd FILL
XFILL_4_CLKBUF1_18 gnd vdd FILL
XFILL_19_7_2 gnd vdd FILL
XFILL_18_NOR3X1_19 gnd vdd FILL
XFILL_4_CLKBUF1_29 gnd vdd FILL
XFILL_18_2_1 gnd vdd FILL
XFILL_0_INVX1_47 gnd vdd FILL
XFILL_1_AND2X2_6 gnd vdd FILL
XFILL_5_INVX8_4 gnd vdd FILL
XFILL_0_INVX1_58 gnd vdd FILL
XFILL_68_DFFSR_208 gnd vdd FILL
XFILL_0_INVX1_69 gnd vdd FILL
XFILL_68_DFFSR_219 gnd vdd FILL
XFILL_18_INVX8_2 gnd vdd FILL
XFILL_46_DFFSR_17 gnd vdd FILL
XFILL_46_DFFSR_28 gnd vdd FILL
XFILL_46_DFFSR_39 gnd vdd FILL
XFILL_31_7 gnd vdd FILL
XFILL_61_5_2 gnd vdd FILL
XFILL_60_0_1 gnd vdd FILL
XFILL_2_NOR2X1_103 gnd vdd FILL
XFILL_24_6 gnd vdd FILL
XFILL_13_OAI21X1_19 gnd vdd FILL
XFILL_86_DFFSR_16 gnd vdd FILL
XFILL_2_NOR2X1_114 gnd vdd FILL
XFILL_2_NOR2X1_125 gnd vdd FILL
XFILL_22_DFFSR_4 gnd vdd FILL
XFILL_86_DFFSR_27 gnd vdd FILL
XFILL_2_NOR2X1_136 gnd vdd FILL
XFILL_2_NOR2X1_147 gnd vdd FILL
XFILL_86_DFFSR_38 gnd vdd FILL
XFILL_17_5 gnd vdd FILL
XFILL_86_DFFSR_49 gnd vdd FILL
XFILL_2_NOR2X1_158 gnd vdd FILL
XFILL_15_DFFSR_16 gnd vdd FILL
XFILL_2_NOR2X1_169 gnd vdd FILL
XFILL_15_DFFSR_27 gnd vdd FILL
XFILL_15_DFFSR_38 gnd vdd FILL
XFILL_15_DFFSR_49 gnd vdd FILL
XFILL_55_DFFSR_15 gnd vdd FILL
XFILL_55_DFFSR_26 gnd vdd FILL
XFILL_55_DFFSR_37 gnd vdd FILL
XFILL_55_DFFSR_48 gnd vdd FILL
XFILL_55_DFFSR_59 gnd vdd FILL
XFILL_53_DFFSR_230 gnd vdd FILL
XFILL_53_DFFSR_241 gnd vdd FILL
XFILL_53_DFFSR_252 gnd vdd FILL
XFILL_53_DFFSR_263 gnd vdd FILL
XFILL_2_MUX2X1_109 gnd vdd FILL
XFILL_53_DFFSR_274 gnd vdd FILL
XFILL_44_DFFSR_8 gnd vdd FILL
XFILL_24_DFFSR_14 gnd vdd FILL
XFILL_7_NOR2X1_203 gnd vdd FILL
XFILL_24_DFFSR_25 gnd vdd FILL
XFILL_80_DFFSR_130 gnd vdd FILL
XFILL_24_DFFSR_36 gnd vdd FILL
XFILL_80_DFFSR_141 gnd vdd FILL
XFILL_57_DFFSR_240 gnd vdd FILL
XFILL_24_DFFSR_47 gnd vdd FILL
XFILL_80_DFFSR_152 gnd vdd FILL
XFILL_24_DFFSR_58 gnd vdd FILL
XFILL_57_DFFSR_251 gnd vdd FILL
XFILL_15_BUFX4_90 gnd vdd FILL
XFILL_57_DFFSR_262 gnd vdd FILL
XFILL_24_DFFSR_69 gnd vdd FILL
XFILL_80_DFFSR_163 gnd vdd FILL
XFILL_80_DFFSR_174 gnd vdd FILL
XFILL_12_CLKBUF1_3 gnd vdd FILL
XFILL_57_DFFSR_273 gnd vdd FILL
XFILL_3_OAI21X1_14 gnd vdd FILL
XFILL_0_DFFSR_200 gnd vdd FILL
XFILL_80_DFFSR_185 gnd vdd FILL
XFILL_0_DFFSR_211 gnd vdd FILL
XFILL_3_OAI21X1_25 gnd vdd FILL
XFILL_80_DFFSR_196 gnd vdd FILL
XFILL_64_DFFSR_13 gnd vdd FILL
XFILL_3_OAI21X1_36 gnd vdd FILL
XFILL_31_DFFSR_209 gnd vdd FILL
XFILL_0_DFFSR_222 gnd vdd FILL
XFILL_64_DFFSR_24 gnd vdd FILL
XFILL_3_OAI21X1_47 gnd vdd FILL
XFILL_64_DFFSR_35 gnd vdd FILL
XFILL_0_DFFSR_233 gnd vdd FILL
XFILL_84_DFFSR_140 gnd vdd FILL
XFILL_64_DFFSR_46 gnd vdd FILL
XFILL_0_DFFSR_244 gnd vdd FILL
XFILL_84_DFFSR_151 gnd vdd FILL
XFILL_0_DFFSR_255 gnd vdd FILL
XFILL_64_DFFSR_57 gnd vdd FILL
XFILL_84_DFFSR_162 gnd vdd FILL
XFILL_64_DFFSR_68 gnd vdd FILL
XFILL_0_DFFSR_266 gnd vdd FILL
XFILL_84_DFFSR_173 gnd vdd FILL
XFILL_64_DFFSR_79 gnd vdd FILL
XFILL_16_CLKBUF1_2 gnd vdd FILL
XFILL_84_DFFSR_184 gnd vdd FILL
XFILL_4_DFFSR_210 gnd vdd FILL
XFILL_84_DFFSR_195 gnd vdd FILL
XFILL_35_DFFSR_208 gnd vdd FILL
XFILL_4_DFFSR_221 gnd vdd FILL
XFILL_52_5_2 gnd vdd FILL
XFILL_35_DFFSR_219 gnd vdd FILL
XFILL_4_DFFSR_232 gnd vdd FILL
XFILL_7_DFFSR_15 gnd vdd FILL
XFILL_4_DFFSR_243 gnd vdd FILL
XFILL_7_DFFSR_26 gnd vdd FILL
XFILL_51_0_1 gnd vdd FILL
XFILL_7_DFFSR_37 gnd vdd FILL
XFILL_4_DFFSR_254 gnd vdd FILL
XFILL_2_NAND2X1_90 gnd vdd FILL
XFILL_33_DFFSR_12 gnd vdd FILL
XFILL_4_DFFSR_265 gnd vdd FILL
XFILL_7_DFFSR_48 gnd vdd FILL
XFILL_33_DFFSR_23 gnd vdd FILL
XFILL_33_DFFSR_34 gnd vdd FILL
XFILL_7_DFFSR_59 gnd vdd FILL
XFILL_33_DFFSR_45 gnd vdd FILL
XFILL_33_DFFSR_56 gnd vdd FILL
XFILL_10_CLKBUF1_10 gnd vdd FILL
XFILL_39_DFFSR_207 gnd vdd FILL
XFILL_10_CLKBUF1_21 gnd vdd FILL
XFILL_62_DFFSR_108 gnd vdd FILL
XFILL_8_DFFSR_220 gnd vdd FILL
XFILL_10_CLKBUF1_32 gnd vdd FILL
XFILL_33_DFFSR_67 gnd vdd FILL
XFILL_62_DFFSR_119 gnd vdd FILL
XFILL_39_DFFSR_218 gnd vdd FILL
XFILL_33_DFFSR_78 gnd vdd FILL
XFILL_8_DFFSR_231 gnd vdd FILL
XFILL_33_DFFSR_89 gnd vdd FILL
XFILL_8_DFFSR_242 gnd vdd FILL
XFILL_39_DFFSR_229 gnd vdd FILL
XFILL_73_DFFSR_11 gnd vdd FILL
XFILL_8_DFFSR_253 gnd vdd FILL
XFILL_8_DFFSR_264 gnd vdd FILL
XFILL_8_DFFSR_275 gnd vdd FILL
XFILL_73_DFFSR_22 gnd vdd FILL
XFILL_73_DFFSR_33 gnd vdd FILL
XFILL_16_MUX2X1_1 gnd vdd FILL
XFILL_73_DFFSR_44 gnd vdd FILL
XFILL_73_DFFSR_55 gnd vdd FILL
XFILL_66_DFFSR_107 gnd vdd FILL
XFILL_73_DFFSR_66 gnd vdd FILL
XFILL_66_DFFSR_118 gnd vdd FILL
XFILL_73_DFFSR_77 gnd vdd FILL
XFILL_66_DFFSR_129 gnd vdd FILL
XFILL_73_DFFSR_88 gnd vdd FILL
XFILL_73_DFFSR_99 gnd vdd FILL
XFILL_9_MUX2X1_19 gnd vdd FILL
XFILL_42_DFFSR_10 gnd vdd FILL
XFILL_6_BUFX4_7 gnd vdd FILL
XFILL_42_DFFSR_21 gnd vdd FILL
XFILL_19_MUX2X1_101 gnd vdd FILL
XFILL_42_DFFSR_32 gnd vdd FILL
XFILL_10_NOR2X1_10 gnd vdd FILL
XFILL_42_DFFSR_43 gnd vdd FILL
XFILL_19_MUX2X1_112 gnd vdd FILL
XFILL_10_NOR2X1_21 gnd vdd FILL
XFILL_1_AOI22X1_4 gnd vdd FILL
XFILL_13_NOR3X1_7 gnd vdd FILL
XFILL_19_MUX2X1_123 gnd vdd FILL
XFILL_13_OAI21X1_7 gnd vdd FILL
XFILL_20_DFFSR_230 gnd vdd FILL
XFILL_42_DFFSR_54 gnd vdd FILL
XFILL_10_NOR2X1_32 gnd vdd FILL
XFILL_10_NOR2X1_43 gnd vdd FILL
XFILL_20_DFFSR_241 gnd vdd FILL
XFILL_42_DFFSR_65 gnd vdd FILL
XFILL_19_MUX2X1_134 gnd vdd FILL
XFILL_42_DFFSR_76 gnd vdd FILL
XFILL_19_MUX2X1_145 gnd vdd FILL
XFILL_10_NOR2X1_54 gnd vdd FILL
XFILL_20_DFFSR_252 gnd vdd FILL
XFILL_19_MUX2X1_156 gnd vdd FILL
XFILL_20_DFFSR_263 gnd vdd FILL
XFILL_10_NOR2X1_65 gnd vdd FILL
XFILL_42_DFFSR_87 gnd vdd FILL
XFILL_20_DFFSR_274 gnd vdd FILL
XFILL_10_NOR2X1_76 gnd vdd FILL
XFILL_42_DFFSR_98 gnd vdd FILL
XFILL_1_INVX1_203 gnd vdd FILL
XFILL_19_MUX2X1_167 gnd vdd FILL
XFILL_59_1_1 gnd vdd FILL
XFILL_82_DFFSR_20 gnd vdd FILL
XFILL_19_MUX2X1_178 gnd vdd FILL
XFILL_1_INVX1_214 gnd vdd FILL
XFILL_10_NOR2X1_87 gnd vdd FILL
XFILL_19_MUX2X1_189 gnd vdd FILL
XFILL_10_NOR2X1_98 gnd vdd FILL
XFILL_82_DFFSR_31 gnd vdd FILL
XFILL_1_INVX1_225 gnd vdd FILL
XFILL_82_DFFSR_42 gnd vdd FILL
XFILL_5_AOI22X1_3 gnd vdd FILL
XFILL_82_DFFSR_53 gnd vdd FILL
XFILL_11_DFFSR_20 gnd vdd FILL
XFILL_24_DFFSR_240 gnd vdd FILL
XFILL_82_DFFSR_64 gnd vdd FILL
XFILL_24_DFFSR_251 gnd vdd FILL
XFILL_11_DFFSR_31 gnd vdd FILL
XFILL_82_DFFSR_75 gnd vdd FILL
XFILL_82_DFFSR_86 gnd vdd FILL
XFILL_24_DFFSR_262 gnd vdd FILL
XFILL_11_DFFSR_42 gnd vdd FILL
XFILL_24_DFFSR_273 gnd vdd FILL
XFILL_5_INVX1_202 gnd vdd FILL
XFILL_11_DFFSR_53 gnd vdd FILL
XFILL_82_DFFSR_97 gnd vdd FILL
XFILL_21_MUX2X1_18 gnd vdd FILL
XFILL_9_NOR2X1_2 gnd vdd FILL
XFILL_5_INVX1_213 gnd vdd FILL
XFILL_11_DFFSR_64 gnd vdd FILL
XFILL_21_MUX2X1_29 gnd vdd FILL
XFILL_11_DFFSR_75 gnd vdd FILL
XFILL_5_INVX1_224 gnd vdd FILL
XFILL_11_DFFSR_86 gnd vdd FILL
XFILL_9_AOI22X1_2 gnd vdd FILL
XFILL_51_DFFSR_140 gnd vdd FILL
XFILL_11_DFFSR_97 gnd vdd FILL
XFILL_51_DFFSR_151 gnd vdd FILL
XFILL_51_DFFSR_30 gnd vdd FILL
XFILL_28_DFFSR_250 gnd vdd FILL
XFILL_2_BUFX2_3 gnd vdd FILL
XFILL_51_DFFSR_162 gnd vdd FILL
XFILL_51_DFFSR_41 gnd vdd FILL
XFILL_28_DFFSR_261 gnd vdd FILL
XFILL_22_NOR3X1_5 gnd vdd FILL
XFILL_43_5_2 gnd vdd FILL
XFILL_28_DFFSR_272 gnd vdd FILL
XFILL_51_DFFSR_173 gnd vdd FILL
XFILL_51_DFFSR_184 gnd vdd FILL
XFILL_51_DFFSR_52 gnd vdd FILL
XFILL_51_DFFSR_63 gnd vdd FILL
XFILL_42_0_1 gnd vdd FILL
XFILL_51_DFFSR_195 gnd vdd FILL
XFILL_51_DFFSR_74 gnd vdd FILL
XFILL_51_DFFSR_85 gnd vdd FILL
XFILL_51_DFFSR_96 gnd vdd FILL
XFILL_55_DFFSR_150 gnd vdd FILL
XFILL_55_DFFSR_161 gnd vdd FILL
XFILL_55_DFFSR_172 gnd vdd FILL
XFILL_55_DFFSR_183 gnd vdd FILL
XFILL_55_DFFSR_194 gnd vdd FILL
XFILL_61_DFFSR_2 gnd vdd FILL
XFILL_20_DFFSR_40 gnd vdd FILL
XFILL_20_DFFSR_51 gnd vdd FILL
XFILL_9_MUX2X1_140 gnd vdd FILL
XFILL_20_DFFSR_62 gnd vdd FILL
XFILL_9_MUX2X1_151 gnd vdd FILL
XFILL_59_DFFSR_160 gnd vdd FILL
XFILL_9_MUX2X1_162 gnd vdd FILL
XFILL_20_DFFSR_73 gnd vdd FILL
XFILL_20_DFFSR_84 gnd vdd FILL
XFILL_9_MUX2X1_173 gnd vdd FILL
XFILL_20_DFFSR_95 gnd vdd FILL
XFILL_9_MUX2X1_184 gnd vdd FILL
XFILL_59_DFFSR_171 gnd vdd FILL
XFILL_5_NOR3X1_6 gnd vdd FILL
XFILL_59_DFFSR_182 gnd vdd FILL
XFILL_59_DFFSR_193 gnd vdd FILL
XFILL_33_DFFSR_107 gnd vdd FILL
XFILL_2_DFFSR_120 gnd vdd FILL
XFILL_2_DFFSR_131 gnd vdd FILL
XFILL_31_NOR3X1_3 gnd vdd FILL
XFILL_33_DFFSR_118 gnd vdd FILL
XFILL_10_NAND2X1_9 gnd vdd FILL
XFILL_2_DFFSR_142 gnd vdd FILL
XFILL_33_DFFSR_129 gnd vdd FILL
XFILL_60_DFFSR_50 gnd vdd FILL
XFILL_2_DFFSR_153 gnd vdd FILL
XFILL_60_DFFSR_61 gnd vdd FILL
XFILL_60_DFFSR_72 gnd vdd FILL
XFILL_2_DFFSR_164 gnd vdd FILL
XFILL_60_DFFSR_83 gnd vdd FILL
XFILL_2_DFFSR_175 gnd vdd FILL
XFILL_2_DFFSR_186 gnd vdd FILL
XFILL_60_DFFSR_94 gnd vdd FILL
XFILL_2_DFFSR_197 gnd vdd FILL
XFILL_37_DFFSR_106 gnd vdd FILL
XFILL_6_DFFSR_130 gnd vdd FILL
XFILL_37_DFFSR_117 gnd vdd FILL
XFILL_3_DFFSR_30 gnd vdd FILL
XFILL_37_DFFSR_128 gnd vdd FILL
XFILL_6_DFFSR_141 gnd vdd FILL
XFILL_6_DFFSR_152 gnd vdd FILL
XFILL_3_DFFSR_41 gnd vdd FILL
XFILL_37_DFFSR_139 gnd vdd FILL
XFILL_10_MUX2X1_50 gnd vdd FILL
XFILL_26_DFFSR_5 gnd vdd FILL
XFILL_11_NAND3X1_15 gnd vdd FILL
XFILL_3_DFFSR_52 gnd vdd FILL
XFILL_11_NAND3X1_26 gnd vdd FILL
XFILL_6_DFFSR_163 gnd vdd FILL
XFILL_10_MUX2X1_61 gnd vdd FILL
XFILL_3_DFFSR_63 gnd vdd FILL
XFILL_6_DFFSR_174 gnd vdd FILL
XFILL_83_DFFSR_6 gnd vdd FILL
XFILL_10_MUX2X1_72 gnd vdd FILL
XFILL_10_MUX2X1_83 gnd vdd FILL
XFILL_3_DFFSR_74 gnd vdd FILL
XFILL_11_NAND3X1_37 gnd vdd FILL
XFILL_6_DFFSR_185 gnd vdd FILL
XFILL_10_MUX2X1_94 gnd vdd FILL
XFILL_3_DFFSR_85 gnd vdd FILL
XFILL_11_NAND3X1_48 gnd vdd FILL
XFILL_6_DFFSR_196 gnd vdd FILL
XFILL_11_NAND3X1_59 gnd vdd FILL
XFILL_3_DFFSR_96 gnd vdd FILL
XFILL_2_INVX2_3 gnd vdd FILL
XFILL_31_CLKBUF1_15 gnd vdd FILL
XFILL_31_CLKBUF1_26 gnd vdd FILL
XFILL_31_CLKBUF1_37 gnd vdd FILL
XFILL_14_MUX2X1_60 gnd vdd FILL
XFILL_14_MUX2X1_71 gnd vdd FILL
XFILL_14_MUX2X1_82 gnd vdd FILL
XFILL_2_NOR3X1_20 gnd vdd FILL
XFILL_14_MUX2X1_93 gnd vdd FILL
XFILL_2_NOR3X1_31 gnd vdd FILL
XFILL_2_NOR3X1_42 gnd vdd FILL
XFILL_83_DFFSR_207 gnd vdd FILL
XFILL_34_5_2 gnd vdd FILL
XFILL_83_DFFSR_218 gnd vdd FILL
XFILL_0_INVX1_1 gnd vdd FILL
XFILL_18_MUX2X1_70 gnd vdd FILL
XFILL_83_DFFSR_229 gnd vdd FILL
XFILL_33_0_1 gnd vdd FILL
XFILL_18_MUX2X1_81 gnd vdd FILL
XFILL_18_MUX2X1_92 gnd vdd FILL
XFILL_22_3 gnd vdd FILL
XFILL_6_NOR3X1_30 gnd vdd FILL
XFILL_6_NOR3X1_41 gnd vdd FILL
XFILL_48_DFFSR_9 gnd vdd FILL
XFILL_6_NOR3X1_52 gnd vdd FILL
XFILL_87_DFFSR_206 gnd vdd FILL
XFILL_15_2 gnd vdd FILL
XFILL_87_DFFSR_217 gnd vdd FILL
XFILL_87_DFFSR_228 gnd vdd FILL
XFILL_22_DFFSR_150 gnd vdd FILL
XFILL_87_DFFSR_239 gnd vdd FILL
XFILL_22_DFFSR_161 gnd vdd FILL
XFILL_22_DFFSR_172 gnd vdd FILL
XFILL_3_INVX1_101 gnd vdd FILL
XFILL_22_DFFSR_183 gnd vdd FILL
XFILL_3_INVX1_112 gnd vdd FILL
XFILL_22_DFFSR_194 gnd vdd FILL
XFILL_3_INVX1_123 gnd vdd FILL
XFILL_3_INVX1_134 gnd vdd FILL
XFILL_1_NAND3X1_10 gnd vdd FILL
XFILL_1_NAND3X1_21 gnd vdd FILL
XFILL_3_INVX1_145 gnd vdd FILL
XFILL_3_INVX1_156 gnd vdd FILL
XFILL_1_NAND3X1_32 gnd vdd FILL
XFILL_1_NAND3X1_43 gnd vdd FILL
XFILL_26_DFFSR_160 gnd vdd FILL
XFILL_3_INVX1_167 gnd vdd FILL
XFILL_5_NAND2X1_12 gnd vdd FILL
XFILL_1_NAND3X1_54 gnd vdd FILL
XFILL_3_INVX1_178 gnd vdd FILL
XFILL_7_INVX1_100 gnd vdd FILL
XFILL_1_NAND3X1_65 gnd vdd FILL
XFILL_3_INVX1_189 gnd vdd FILL
XFILL_5_NAND2X1_23 gnd vdd FILL
XFILL_26_DFFSR_171 gnd vdd FILL
XFILL_1_NAND3X1_76 gnd vdd FILL
XFILL_7_INVX1_111 gnd vdd FILL
XFILL_26_DFFSR_182 gnd vdd FILL
XFILL_1_NAND3X1_87 gnd vdd FILL
XFILL_26_DFFSR_193 gnd vdd FILL
XFILL_5_NAND2X1_34 gnd vdd FILL
XFILL_7_INVX1_122 gnd vdd FILL
XFILL_5_NAND2X1_45 gnd vdd FILL
XFILL_1_NAND3X1_98 gnd vdd FILL
XFILL_7_INVX1_133 gnd vdd FILL
XFILL_5_NAND2X1_56 gnd vdd FILL
XFILL_7_INVX1_144 gnd vdd FILL
XFILL_5_NAND2X1_67 gnd vdd FILL
XFILL_7_INVX1_155 gnd vdd FILL
XFILL_5_NAND2X1_78 gnd vdd FILL
XINVX1_180 INVX1_180/A gnd INVX1_180/Y vdd INVX1
XFILL_5_NAND2X1_89 gnd vdd FILL
XFILL_7_INVX1_166 gnd vdd FILL
XINVX1_191 INVX1_191/A gnd INVX1_191/Y vdd INVX1
XFILL_7_INVX1_177 gnd vdd FILL
XFILL_7_INVX1_188 gnd vdd FILL
XFILL_7_INVX1_199 gnd vdd FILL
XFILL_22_NOR3X1_50 gnd vdd FILL
XFILL_1_OAI22X1_7 gnd vdd FILL
XFILL_72_DFFSR_250 gnd vdd FILL
XFILL_72_DFFSR_261 gnd vdd FILL
XFILL_72_DFFSR_272 gnd vdd FILL
XFILL_5_OAI22X1_6 gnd vdd FILL
XFILL_11_NOR2X1_105 gnd vdd FILL
XFILL_11_NOR2X1_116 gnd vdd FILL
XFILL_11_NOR2X1_127 gnd vdd FILL
XFILL_11_NOR2X1_138 gnd vdd FILL
XFILL_5_AOI22X1_10 gnd vdd FILL
XFILL_76_DFFSR_260 gnd vdd FILL
XFILL_25_5_2 gnd vdd FILL
XFILL_76_DFFSR_271 gnd vdd FILL
XFILL_11_NOR2X1_149 gnd vdd FILL
XFILL_31_CLKBUF1_1 gnd vdd FILL
XFILL_0_5_2 gnd vdd FILL
XFILL_24_0_1 gnd vdd FILL
XFILL_50_DFFSR_207 gnd vdd FILL
XFILL_9_AOI21X1_12 gnd vdd FILL
XFILL_9_OAI22X1_5 gnd vdd FILL
XFILL_50_DFFSR_218 gnd vdd FILL
XFILL_9_AOI21X1_23 gnd vdd FILL
XFILL_50_DFFSR_229 gnd vdd FILL
XFILL_9_AOI21X1_34 gnd vdd FILL
XFILL_9_AOI21X1_45 gnd vdd FILL
XFILL_9_AOI21X1_56 gnd vdd FILL
XFILL_9_AOI21X1_67 gnd vdd FILL
XFILL_19_OAI22X1_14 gnd vdd FILL
XFILL_20_CLKBUF1_11 gnd vdd FILL
XFILL_9_AOI21X1_78 gnd vdd FILL
XFILL_19_OAI22X1_25 gnd vdd FILL
XFILL_19_OAI22X1_36 gnd vdd FILL
XFILL_54_DFFSR_206 gnd vdd FILL
XFILL_20_CLKBUF1_22 gnd vdd FILL
XFILL_19_OAI22X1_47 gnd vdd FILL
XFILL_54_DFFSR_217 gnd vdd FILL
XFILL_20_CLKBUF1_33 gnd vdd FILL
XFILL_54_DFFSR_228 gnd vdd FILL
XFILL_54_DFFSR_239 gnd vdd FILL
XFILL_3_CLKBUF1_15 gnd vdd FILL
XFILL_3_CLKBUF1_26 gnd vdd FILL
XFILL_3_CLKBUF1_37 gnd vdd FILL
XFILL_81_DFFSR_106 gnd vdd FILL
XFILL_58_DFFSR_205 gnd vdd FILL
XFILL_58_DFFSR_216 gnd vdd FILL
XFILL_81_DFFSR_117 gnd vdd FILL
XFILL_58_DFFSR_227 gnd vdd FILL
XFILL_81_DFFSR_128 gnd vdd FILL
XFILL_81_DFFSR_139 gnd vdd FILL
XFILL_58_DFFSR_238 gnd vdd FILL
XFILL_6_BUFX2_4 gnd vdd FILL
XFILL_58_DFFSR_249 gnd vdd FILL
XFILL_85_DFFSR_105 gnd vdd FILL
XFILL_1_NOR2X1_100 gnd vdd FILL
XFILL_1_DFFSR_209 gnd vdd FILL
XFILL_1_NOR2X1_111 gnd vdd FILL
XFILL_12_OAI21X1_16 gnd vdd FILL
XFILL_85_DFFSR_116 gnd vdd FILL
XFILL_12_OAI21X1_27 gnd vdd FILL
XFILL_85_DFFSR_127 gnd vdd FILL
XFILL_1_NOR2X1_122 gnd vdd FILL
XFILL_85_DFFSR_138 gnd vdd FILL
XFILL_1_NOR2X1_133 gnd vdd FILL
XFILL_8_6_2 gnd vdd FILL
XFILL_85_DFFSR_149 gnd vdd FILL
XFILL_1_NOR2X1_144 gnd vdd FILL
XFILL_12_OAI21X1_38 gnd vdd FILL
XFILL_12_OAI21X1_49 gnd vdd FILL
XFILL_1_NOR2X1_155 gnd vdd FILL
XFILL_7_1_1 gnd vdd FILL
XFILL_1_NOR2X1_166 gnd vdd FILL
XFILL_65_DFFSR_3 gnd vdd FILL
XFILL_1_NOR2X1_177 gnd vdd FILL
XFILL_8_BUFX4_12 gnd vdd FILL
XFILL_5_DFFSR_208 gnd vdd FILL
XFILL_1_NOR2X1_188 gnd vdd FILL
XFILL_5_DFFSR_219 gnd vdd FILL
XFILL_8_BUFX4_23 gnd vdd FILL
XFILL_1_NOR2X1_199 gnd vdd FILL
XFILL_2_NAND3X1_8 gnd vdd FILL
XFILL_8_BUFX4_34 gnd vdd FILL
XFILL_8_BUFX4_45 gnd vdd FILL
XFILL_8_BUFX4_56 gnd vdd FILL
XFILL_9_OAI22X1_20 gnd vdd FILL
XFILL_11_NAND2X1_70 gnd vdd FILL
XFILL_8_BUFX4_67 gnd vdd FILL
XFILL_11_NAND2X1_81 gnd vdd FILL
XFILL_9_OAI22X1_31 gnd vdd FILL
XFILL_8_BUFX4_78 gnd vdd FILL
XFILL_11_NAND2X1_92 gnd vdd FILL
XFILL_9_OAI22X1_42 gnd vdd FILL
XFILL_8_BUFX4_89 gnd vdd FILL
XFILL_9_DFFSR_207 gnd vdd FILL
XFILL_6_NAND3X1_7 gnd vdd FILL
XFILL_9_DFFSR_218 gnd vdd FILL
XFILL_9_DFFSR_229 gnd vdd FILL
XFILL_16_5_2 gnd vdd FILL
XFILL_15_0_1 gnd vdd FILL
XFILL_43_DFFSR_260 gnd vdd FILL
XNAND3X1_100 INVX2_5/Y OAI21X1_43/Y NAND3X1_36/C gnd NAND3X1_39/B vdd NAND3X1
XFILL_43_DFFSR_271 gnd vdd FILL
XFILL_1_MUX2X1_106 gnd vdd FILL
XNAND3X1_111 NOR3X1_9/A DFFSR_199/D AND2X2_3/B gnd NOR3X1_39/C vdd NAND3X1
XFILL_1_MUX2X1_117 gnd vdd FILL
XNAND3X1_122 INVX2_2/A AND2X2_5/B NAND3X1_2/C gnd OAI22X1_1/D vdd NAND3X1
XFILL_1_MUX2X1_128 gnd vdd FILL
XFILL_6_NOR2X1_200 gnd vdd FILL
XFILL_1_MUX2X1_139 gnd vdd FILL
XFILL_87_DFFSR_7 gnd vdd FILL
XFILL_70_DFFSR_160 gnd vdd FILL
XFILL_47_DFFSR_270 gnd vdd FILL
XFILL_70_DFFSR_171 gnd vdd FILL
XFILL_2_OAI21X1_11 gnd vdd FILL
XFILL_6_INVX2_4 gnd vdd FILL
XFILL_70_DFFSR_182 gnd vdd FILL
XFILL_52_DFFSR_19 gnd vdd FILL
XFILL_70_DFFSR_193 gnd vdd FILL
XFILL_2_OAI21X1_22 gnd vdd FILL
XFILL_21_DFFSR_206 gnd vdd FILL
XFILL_2_OAI21X1_33 gnd vdd FILL
XFILL_21_DFFSR_217 gnd vdd FILL
XFILL_2_OAI21X1_44 gnd vdd FILL
XFILL_11_NOR2X1_19 gnd vdd FILL
XFILL_21_DFFSR_228 gnd vdd FILL
XFILL_21_DFFSR_239 gnd vdd FILL
XFILL_74_DFFSR_170 gnd vdd FILL
XFILL_74_DFFSR_181 gnd vdd FILL
XFILL_74_DFFSR_192 gnd vdd FILL
XFILL_25_DFFSR_205 gnd vdd FILL
XFILL_15_AOI21X1_70 gnd vdd FILL
XFILL_25_DFFSR_216 gnd vdd FILL
XFILL_15_AOI21X1_81 gnd vdd FILL
XFILL_4_INVX1_2 gnd vdd FILL
XFILL_25_DFFSR_227 gnd vdd FILL
XFILL_25_DFFSR_238 gnd vdd FILL
XFILL_21_DFFSR_18 gnd vdd FILL
XFILL_12_BUFX4_50 gnd vdd FILL
XFILL_25_DFFSR_249 gnd vdd FILL
XFILL_21_DFFSR_29 gnd vdd FILL
XFILL_12_BUFX4_61 gnd vdd FILL
XFILL_12_BUFX4_72 gnd vdd FILL
XFILL_78_DFFSR_180 gnd vdd FILL
XFILL_12_BUFX4_83 gnd vdd FILL
XFILL_78_DFFSR_191 gnd vdd FILL
XFILL_52_DFFSR_105 gnd vdd FILL
XFILL_29_DFFSR_204 gnd vdd FILL
XFILL_12_BUFX4_94 gnd vdd FILL
XFILL_29_DFFSR_215 gnd vdd FILL
XFILL_52_DFFSR_116 gnd vdd FILL
XFILL_52_DFFSR_127 gnd vdd FILL
XFILL_29_DFFSR_226 gnd vdd FILL
XFILL_52_DFFSR_138 gnd vdd FILL
XFILL_52_DFFSR_149 gnd vdd FILL
XFILL_29_DFFSR_237 gnd vdd FILL
XFILL_61_DFFSR_17 gnd vdd FILL
XFILL_29_DFFSR_248 gnd vdd FILL
XFILL_61_DFFSR_28 gnd vdd FILL
XFILL_61_DFFSR_39 gnd vdd FILL
XFILL_29_DFFSR_259 gnd vdd FILL
XFILL_66_4_2 gnd vdd FILL
XFILL_56_DFFSR_104 gnd vdd FILL
XFILL_56_DFFSR_115 gnd vdd FILL
XFILL_56_DFFSR_126 gnd vdd FILL
XFILL_56_DFFSR_137 gnd vdd FILL
XFILL_56_DFFSR_148 gnd vdd FILL
XFILL_56_DFFSR_159 gnd vdd FILL
XFILL_4_DFFSR_19 gnd vdd FILL
XFILL_30_DFFSR_16 gnd vdd FILL
XFILL_30_DFFSR_27 gnd vdd FILL
XFILL_30_DFFSR_38 gnd vdd FILL
XFILL_30_DFFSR_49 gnd vdd FILL
XFILL_6_INVX1_40 gnd vdd FILL
XFILL_6_INVX1_51 gnd vdd FILL
XFILL_18_MUX2X1_120 gnd vdd FILL
XFILL_6_INVX1_62 gnd vdd FILL
XFILL_18_MUX2X1_131 gnd vdd FILL
XFILL_18_MUX2X1_142 gnd vdd FILL
XFILL_6_INVX1_73 gnd vdd FILL
XFILL_18_MUX2X1_153 gnd vdd FILL
XFILL_6_INVX1_84 gnd vdd FILL
XFILL_10_DFFSR_260 gnd vdd FILL
XFILL_10_DFFSR_271 gnd vdd FILL
XFILL_18_MUX2X1_164 gnd vdd FILL
XFILL_6_INVX1_95 gnd vdd FILL
XFILL_70_DFFSR_15 gnd vdd FILL
XFILL_3_DFFSR_107 gnd vdd FILL
XFILL_18_MUX2X1_175 gnd vdd FILL
XFILL_70_DFFSR_26 gnd vdd FILL
XFILL_3_DFFSR_118 gnd vdd FILL
XFILL_70_DFFSR_37 gnd vdd FILL
XFILL_18_MUX2X1_186 gnd vdd FILL
XFILL_3_DFFSR_129 gnd vdd FILL
XFILL_70_DFFSR_48 gnd vdd FILL
XFILL_13_MUX2X1_5 gnd vdd FILL
XFILL_70_DFFSR_59 gnd vdd FILL
XFILL_7_DFFSR_106 gnd vdd FILL
XFILL_14_DFFSR_270 gnd vdd FILL
XDFFSR_120 INVX1_182/A CLKBUF1_31/Y DFFSR_64/R vdd DFFSR_120/D gnd vdd DFFSR
XDFFSR_131 INVX1_167/A DFFSR_55/CLK DFFSR_58/R vdd DFFSR_131/D gnd vdd DFFSR
XFILL_7_DFFSR_117 gnd vdd FILL
XFILL_11_MUX2X1_15 gnd vdd FILL
XDFFSR_142 DFFSR_142/Q CLKBUF1_1/Y DFFSR_58/R vdd DFFSR_142/D gnd vdd DFFSR
XFILL_7_DFFSR_128 gnd vdd FILL
XFILL_11_MUX2X1_26 gnd vdd FILL
XDFFSR_153 INVX1_151/A DFFSR_78/CLK DFFSR_78/R vdd DFFSR_153/D gnd vdd DFFSR
XFILL_11_MUX2X1_37 gnd vdd FILL
XFILL_7_DFFSR_139 gnd vdd FILL
XFILL_4_BUFX4_60 gnd vdd FILL
XFILL_2_AOI21X1_2 gnd vdd FILL
XFILL_11_MUX2X1_48 gnd vdd FILL
XDFFSR_164 INVX1_149/A DFFSR_70/CLK BUFX4_55/Y vdd DFFSR_164/D gnd vdd DFFSR
XDFFSR_175 INVX1_13/A DFFSR_72/CLK BUFX4_55/Y vdd DFFSR_175/D gnd vdd DFFSR
XFILL_4_BUFX4_71 gnd vdd FILL
XBUFX4_5 BUFX4_8/A gnd BUFX4_5/Y vdd BUFX4
XFILL_11_MUX2X1_59 gnd vdd FILL
XFILL_4_BUFX4_82 gnd vdd FILL
XFILL_4_BUFX4_93 gnd vdd FILL
XDFFSR_186 INVX1_112/A DFFSR_70/CLK BUFX4_55/Y vdd DFFSR_186/D gnd vdd DFFSR
XDFFSR_197 INVX1_97/A CLKBUF1_7/Y BUFX4_13/Y vdd MUX2X1_84/Y gnd vdd DFFSR
XFILL_41_DFFSR_170 gnd vdd FILL
XFILL_15_MUX2X1_14 gnd vdd FILL
XFILL_41_DFFSR_181 gnd vdd FILL
XFILL_41_DFFSR_192 gnd vdd FILL
XFILL_15_MUX2X1_25 gnd vdd FILL
XFILL_15_MUX2X1_36 gnd vdd FILL
XFILL_15_MUX2X1_47 gnd vdd FILL
XFILL_6_AOI21X1_1 gnd vdd FILL
XFILL_15_MUX2X1_58 gnd vdd FILL
XFILL_15_MUX2X1_69 gnd vdd FILL
XFILL_3_NOR3X1_18 gnd vdd FILL
XFILL_22_MUX2X1_3 gnd vdd FILL
XFILL_3_NOR3X1_29 gnd vdd FILL
XFILL_45_DFFSR_180 gnd vdd FILL
XFILL_19_MUX2X1_13 gnd vdd FILL
XFILL_45_DFFSR_191 gnd vdd FILL
XFILL_19_MUX2X1_24 gnd vdd FILL
XFILL_19_MUX2X1_35 gnd vdd FILL
XFILL_19_MUX2X1_46 gnd vdd FILL
XFILL_6_NOR2X1_6 gnd vdd FILL
XFILL_57_4_2 gnd vdd FILL
XFILL_19_MUX2X1_57 gnd vdd FILL
XFILL_19_MUX2X1_68 gnd vdd FILL
XNOR3X1_20 NOR3X1_20/A NOR3X1_20/B NOR3X1_20/C gnd NOR3X1_20/Y vdd NOR3X1
XFILL_19_MUX2X1_79 gnd vdd FILL
XFILL_7_NOR3X1_17 gnd vdd FILL
XFILL_8_MUX2X1_170 gnd vdd FILL
XNOR3X1_31 NOR3X1_31/A NOR3X1_31/B NOR3X1_31/C gnd NOR3X1_31/Y vdd NOR3X1
XFILL_7_NOR3X1_28 gnd vdd FILL
XNOR3X1_42 NOR3X1_42/A NOR3X1_42/B NOR3X1_42/C gnd NOR3X1_42/Y vdd NOR3X1
XFILL_8_MUX2X1_181 gnd vdd FILL
XFILL_7_NOR3X1_39 gnd vdd FILL
XFILL_23_DFFSR_104 gnd vdd FILL
XFILL_49_DFFSR_190 gnd vdd FILL
XFILL_8_MUX2X1_192 gnd vdd FILL
XFILL_23_DFFSR_115 gnd vdd FILL
XFILL_23_DFFSR_126 gnd vdd FILL
XFILL_23_DFFSR_137 gnd vdd FILL
XFILL_23_DFFSR_148 gnd vdd FILL
XFILL_23_DFFSR_159 gnd vdd FILL
XFILL_5_MUX2X1_4 gnd vdd FILL
XFILL_27_DFFSR_103 gnd vdd FILL
XFILL_27_DFFSR_114 gnd vdd FILL
XFILL_27_DFFSR_125 gnd vdd FILL
XFILL_27_DFFSR_136 gnd vdd FILL
XFILL_40_3_2 gnd vdd FILL
XFILL_31_DFFSR_6 gnd vdd FILL
XFILL_10_NAND3X1_12 gnd vdd FILL
XFILL_27_DFFSR_147 gnd vdd FILL
XFILL_27_DFFSR_158 gnd vdd FILL
XFILL_10_NAND3X1_23 gnd vdd FILL
XFILL_27_DFFSR_169 gnd vdd FILL
XFILL_10_NAND3X1_34 gnd vdd FILL
XFILL_10_NAND3X1_45 gnd vdd FILL
XFILL_69_DFFSR_4 gnd vdd FILL
XFILL_10_NAND3X1_56 gnd vdd FILL
XFILL_30_CLKBUF1_12 gnd vdd FILL
XFILL_10_NAND3X1_67 gnd vdd FILL
XFILL_10_NAND3X1_78 gnd vdd FILL
XFILL_30_CLKBUF1_23 gnd vdd FILL
XFILL_30_CLKBUF1_34 gnd vdd FILL
XFILL_8_OR2X2_1 gnd vdd FILL
XFILL_10_NAND3X1_89 gnd vdd FILL
XFILL_39_DFFSR_60 gnd vdd FILL
XFILL_39_DFFSR_71 gnd vdd FILL
XFILL_39_DFFSR_82 gnd vdd FILL
XFILL_23_NOR3X1_15 gnd vdd FILL
XFILL_39_DFFSR_93 gnd vdd FILL
XFILL_23_NOR3X1_26 gnd vdd FILL
XFILL_23_NOR3X1_37 gnd vdd FILL
XFILL_23_NOR3X1_48 gnd vdd FILL
XFILL_73_DFFSR_204 gnd vdd FILL
XFILL_73_DFFSR_215 gnd vdd FILL
XFILL_0_DFFSR_12 gnd vdd FILL
XFILL_73_DFFSR_226 gnd vdd FILL
XFILL_0_DFFSR_23 gnd vdd FILL
XFILL_73_DFFSR_237 gnd vdd FILL
XFILL_79_DFFSR_70 gnd vdd FILL
XFILL_0_DFFSR_34 gnd vdd FILL
XFILL_73_DFFSR_248 gnd vdd FILL
XFILL_79_DFFSR_81 gnd vdd FILL
XFILL_0_DFFSR_45 gnd vdd FILL
XFILL_27_NOR3X1_14 gnd vdd FILL
XFILL_0_DFFSR_56 gnd vdd FILL
XFILL_73_DFFSR_259 gnd vdd FILL
XFILL_79_DFFSR_92 gnd vdd FILL
XFILL_27_NOR3X1_25 gnd vdd FILL
XFILL_0_DFFSR_67 gnd vdd FILL
XFILL_27_NOR3X1_36 gnd vdd FILL
XFILL_0_DFFSR_78 gnd vdd FILL
XFILL_0_DFFSR_89 gnd vdd FILL
XFILL_27_NOR3X1_47 gnd vdd FILL
XFILL_77_DFFSR_203 gnd vdd FILL
XFILL_77_DFFSR_214 gnd vdd FILL
XFILL_77_DFFSR_225 gnd vdd FILL
XFILL_1_OAI22X1_19 gnd vdd FILL
XFILL_77_DFFSR_236 gnd vdd FILL
XFILL_77_DFFSR_247 gnd vdd FILL
XFILL_1_CLKBUF1_1 gnd vdd FILL
XFILL_77_DFFSR_258 gnd vdd FILL
XFILL_12_DFFSR_180 gnd vdd FILL
XFILL_77_DFFSR_269 gnd vdd FILL
XFILL_48_4_2 gnd vdd FILL
XFILL_12_DFFSR_191 gnd vdd FILL
XFILL_48_DFFSR_80 gnd vdd FILL
XFILL_48_DFFSR_91 gnd vdd FILL
XFILL_0_NAND3X1_40 gnd vdd FILL
XFILL_0_NAND3X1_51 gnd vdd FILL
XFILL_0_NAND3X1_62 gnd vdd FILL
XFILL_4_NAND2X1_20 gnd vdd FILL
XFILL_0_NAND3X1_73 gnd vdd FILL
XFILL_4_NAND2X1_31 gnd vdd FILL
XFILL_0_NAND3X1_84 gnd vdd FILL
XFILL_16_DFFSR_190 gnd vdd FILL
XFILL_0_NAND3X1_95 gnd vdd FILL
XFILL_4_NAND2X1_42 gnd vdd FILL
XFILL_4_NAND2X1_53 gnd vdd FILL
XFILL_4_NAND2X1_64 gnd vdd FILL
XFILL_4_NAND2X1_75 gnd vdd FILL
XFILL_4_NAND2X1_86 gnd vdd FILL
XFILL_17_DFFSR_90 gnd vdd FILL
XFILL_31_3_2 gnd vdd FILL
XFILL_12_CLKBUF1_17 gnd vdd FILL
XFILL_12_CLKBUF1_28 gnd vdd FILL
XFILL_12_CLKBUF1_39 gnd vdd FILL
XFILL_10_NOR2X1_102 gnd vdd FILL
XFILL_10_NOR2X1_113 gnd vdd FILL
XFILL_10_NOR2X1_124 gnd vdd FILL
XFILL_10_NOR2X1_135 gnd vdd FILL
XFILL_10_NOR2X1_146 gnd vdd FILL
XFILL_10_NOR2X1_157 gnd vdd FILL
XFILL_10_NOR2X1_168 gnd vdd FILL
XFILL_10_NOR2X1_179 gnd vdd FILL
XFILL_40_DFFSR_204 gnd vdd FILL
XFILL_40_DFFSR_215 gnd vdd FILL
XFILL_8_AOI21X1_20 gnd vdd FILL
XFILL_2_OAI21X1_5 gnd vdd FILL
XFILL_8_AOI21X1_31 gnd vdd FILL
XFILL_40_DFFSR_226 gnd vdd FILL
XFILL_40_DFFSR_237 gnd vdd FILL
XFILL_8_AOI21X1_42 gnd vdd FILL
XFILL_40_DFFSR_248 gnd vdd FILL
XFILL_18_OAI22X1_11 gnd vdd FILL
XFILL_8_AOI21X1_53 gnd vdd FILL
XFILL_40_DFFSR_259 gnd vdd FILL
XNAND3X1_8 NAND3X1_8/A NAND3X1_8/B NAND3X1_8/C gnd NOR2X1_97/A vdd NAND3X1
XFILL_8_AOI21X1_64 gnd vdd FILL
XFILL_8_AOI21X1_75 gnd vdd FILL
XFILL_18_OAI22X1_22 gnd vdd FILL
XFILL_18_OAI22X1_33 gnd vdd FILL
XFILL_18_OAI22X1_44 gnd vdd FILL
XFILL_44_DFFSR_203 gnd vdd FILL
XFILL_44_DFFSR_214 gnd vdd FILL
XFILL_6_OAI21X1_4 gnd vdd FILL
XFILL_44_DFFSR_225 gnd vdd FILL
XFILL_39_4_2 gnd vdd FILL
XFILL_3_NOR2X1_40 gnd vdd FILL
XFILL_3_NOR2X1_51 gnd vdd FILL
XFILL_44_DFFSR_236 gnd vdd FILL
XFILL_3_NOR2X1_62 gnd vdd FILL
XFILL_44_DFFSR_247 gnd vdd FILL
XFILL_2_CLKBUF1_12 gnd vdd FILL
XFILL_44_DFFSR_258 gnd vdd FILL
XFILL_3_NOR2X1_73 gnd vdd FILL
XFILL_44_DFFSR_269 gnd vdd FILL
XFILL_2_CLKBUF1_23 gnd vdd FILL
XFILL_13_BUFX4_17 gnd vdd FILL
XFILL_13_BUFX4_28 gnd vdd FILL
XFILL_2_CLKBUF1_34 gnd vdd FILL
XFILL_3_NOR2X1_84 gnd vdd FILL
XFILL_3_NOR2X1_95 gnd vdd FILL
XFILL_71_DFFSR_103 gnd vdd FILL
XFILL_13_BUFX4_39 gnd vdd FILL
XFILL_48_DFFSR_202 gnd vdd FILL
XFILL_10_MUX2X1_108 gnd vdd FILL
XFILL_48_DFFSR_213 gnd vdd FILL
XFILL_71_DFFSR_114 gnd vdd FILL
XFILL_10_MUX2X1_119 gnd vdd FILL
XFILL_48_DFFSR_224 gnd vdd FILL
XFILL_71_DFFSR_125 gnd vdd FILL
XFILL_71_DFFSR_136 gnd vdd FILL
XFILL_48_DFFSR_235 gnd vdd FILL
XFILL_11_OAI22X1_1 gnd vdd FILL
XFILL_71_DFFSR_147 gnd vdd FILL
XFILL_7_NOR2X1_50 gnd vdd FILL
XFILL_71_DFFSR_158 gnd vdd FILL
XFILL_7_NOR2X1_61 gnd vdd FILL
XFILL_48_DFFSR_246 gnd vdd FILL
XFILL_48_DFFSR_257 gnd vdd FILL
XFILL_7_NOR2X1_72 gnd vdd FILL
XFILL_48_DFFSR_268 gnd vdd FILL
XFILL_71_DFFSR_169 gnd vdd FILL
XFILL_7_NOR2X1_83 gnd vdd FILL
XFILL_75_DFFSR_102 gnd vdd FILL
XFILL_7_NOR2X1_94 gnd vdd FILL
XFILL_75_DFFSR_113 gnd vdd FILL
XFILL_11_OAI21X1_13 gnd vdd FILL
XFILL_75_DFFSR_124 gnd vdd FILL
XFILL_50_6_0 gnd vdd FILL
XFILL_11_OAI21X1_24 gnd vdd FILL
XFILL_0_DFFSR_5 gnd vdd FILL
XFILL_75_DFFSR_135 gnd vdd FILL
XFILL_11_OAI21X1_35 gnd vdd FILL
XFILL_22_3_2 gnd vdd FILL
XFILL_0_NOR2X1_130 gnd vdd FILL
XFILL_75_DFFSR_146 gnd vdd FILL
XFILL_0_NOR2X1_141 gnd vdd FILL
XFILL_13_DFFSR_3 gnd vdd FILL
XFILL_75_DFFSR_157 gnd vdd FILL
XFILL_11_OAI21X1_46 gnd vdd FILL
XFILL_0_NOR2X1_152 gnd vdd FILL
XFILL_75_DFFSR_168 gnd vdd FILL
XFILL_0_NOR2X1_163 gnd vdd FILL
XFILL_70_DFFSR_4 gnd vdd FILL
XFILL_75_DFFSR_179 gnd vdd FILL
XFILL_0_NOR2X1_174 gnd vdd FILL
XFILL_79_DFFSR_101 gnd vdd FILL
XFILL_0_NOR2X1_185 gnd vdd FILL
XFILL_79_DFFSR_112 gnd vdd FILL
XFILL_0_NOR2X1_196 gnd vdd FILL
XFILL_79_DFFSR_123 gnd vdd FILL
XFILL_79_DFFSR_134 gnd vdd FILL
XFILL_79_DFFSR_145 gnd vdd FILL
XFILL_79_DFFSR_156 gnd vdd FILL
XFILL_7_INVX1_18 gnd vdd FILL
XFILL_79_DFFSR_167 gnd vdd FILL
XFILL_7_INVX1_29 gnd vdd FILL
XFILL_79_DFFSR_178 gnd vdd FILL
XFILL_8_OAI22X1_50 gnd vdd FILL
XFILL_79_DFFSR_189 gnd vdd FILL
XBUFX2_2 BUFX2_2/A gnd dout[2] vdd BUFX2
XFILL_0_MUX2X1_103 gnd vdd FILL
XFILL_0_MUX2X1_114 gnd vdd FILL
XFILL_0_MUX2X1_125 gnd vdd FILL
XFILL_3_NAND2X1_6 gnd vdd FILL
XFILL_0_MUX2X1_136 gnd vdd FILL
XFILL_35_DFFSR_7 gnd vdd FILL
XFILL_5_BUFX4_16 gnd vdd FILL
XFILL_0_MUX2X1_147 gnd vdd FILL
XFILL_5_BUFX4_27 gnd vdd FILL
XFILL_0_MUX2X1_158 gnd vdd FILL
XFILL_0_MUX2X1_169 gnd vdd FILL
XFILL_5_BUFX4_38 gnd vdd FILL
XFILL_5_BUFX4_49 gnd vdd FILL
XFILL_58_7_0 gnd vdd FILL
XFILL_60_DFFSR_190 gnd vdd FILL
XFILL_5_4_2 gnd vdd FILL
XFILL_7_NAND2X1_5 gnd vdd FILL
XFILL_1_OAI21X1_30 gnd vdd FILL
XFILL_11_DFFSR_203 gnd vdd FILL
XFILL_1_OAI21X1_41 gnd vdd FILL
XFILL_11_DFFSR_214 gnd vdd FILL
XFILL_11_DFFSR_225 gnd vdd FILL
XFILL_11_DFFSR_236 gnd vdd FILL
XFILL_3_MUX2X1_80 gnd vdd FILL
XFILL_11_DFFSR_247 gnd vdd FILL
XFILL_3_MUX2X1_91 gnd vdd FILL
XFILL_11_DFFSR_258 gnd vdd FILL
XFILL_11_DFFSR_269 gnd vdd FILL
XFILL_15_DFFSR_202 gnd vdd FILL
XFILL_15_DFFSR_213 gnd vdd FILL
XFILL_12_NAND3X1_2 gnd vdd FILL
XFILL_15_DFFSR_224 gnd vdd FILL
XFILL_15_DFFSR_235 gnd vdd FILL
XFILL_15_DFFSR_246 gnd vdd FILL
XFILL_7_MUX2X1_90 gnd vdd FILL
XFILL_15_DFFSR_257 gnd vdd FILL
XFILL_15_DFFSR_268 gnd vdd FILL
XFILL_41_6_0 gnd vdd FILL
XFILL_13_3_2 gnd vdd FILL
XFILL_42_DFFSR_102 gnd vdd FILL
XFILL_19_DFFSR_201 gnd vdd FILL
XFILL_12_AND2X2_4 gnd vdd FILL
XFILL_19_DFFSR_212 gnd vdd FILL
XFILL_42_DFFSR_113 gnd vdd FILL
XFILL_42_DFFSR_124 gnd vdd FILL
XFILL_19_DFFSR_223 gnd vdd FILL
XFILL_19_DFFSR_234 gnd vdd FILL
XFILL_42_DFFSR_135 gnd vdd FILL
XINVX2_2 INVX2_2/A gnd INVX2_2/Y vdd INVX2
XFILL_42_DFFSR_146 gnd vdd FILL
XFILL_42_DFFSR_157 gnd vdd FILL
XFILL_19_DFFSR_245 gnd vdd FILL
XFILL_19_DFFSR_256 gnd vdd FILL
XFILL_19_DFFSR_267 gnd vdd FILL
XFILL_42_DFFSR_168 gnd vdd FILL
XFILL_42_DFFSR_179 gnd vdd FILL
XFILL_46_DFFSR_101 gnd vdd FILL
XFILL_46_DFFSR_112 gnd vdd FILL
XAOI21X1_2 BUFX4_72/Y AOI21X1_3/B AOI21X1_2/C gnd DFFSR_150/D vdd AOI21X1
XFILL_3_NAND3X1_17 gnd vdd FILL
XFILL_46_DFFSR_123 gnd vdd FILL
XFILL_46_DFFSR_134 gnd vdd FILL
XFILL_3_NAND3X1_28 gnd vdd FILL
XFILL_46_DFFSR_145 gnd vdd FILL
XFILL_3_NAND3X1_39 gnd vdd FILL
XFILL_46_DFFSR_156 gnd vdd FILL
XFILL_46_DFFSR_167 gnd vdd FILL
XFILL_7_NAND2X1_19 gnd vdd FILL
XFILL_46_DFFSR_178 gnd vdd FILL
XFILL_46_DFFSR_189 gnd vdd FILL
XMUX2X1_160 BUFX4_99/Y INVX1_204/Y NOR2X1_156/Y gnd DFFSR_88/D vdd MUX2X1
XMUX2X1_171 BUFX4_67/Y INVX1_216/Y NOR2X1_165/Y gnd DFFSR_69/D vdd MUX2X1
XMUX2X1_182 BUFX4_98/Y INVX1_227/Y NOR2X1_167/Y gnd DFFSR_62/D vdd MUX2X1
XFILL_12_AOI22X1_7 gnd vdd FILL
XFILL_17_MUX2X1_150 gnd vdd FILL
XMUX2X1_193 MUX2X1_9/A INVX1_14/Y MUX2X1_3/S gnd DFFSR_47/D vdd MUX2X1
XFILL_17_MUX2X1_161 gnd vdd FILL
XFILL_5_5 gnd vdd FILL
XFILL_17_MUX2X1_172 gnd vdd FILL
XFILL_17_MUX2X1_183 gnd vdd FILL
XFILL_17_MUX2X1_194 gnd vdd FILL
XFILL_49_7_0 gnd vdd FILL
XFILL_16_AOI22X1_6 gnd vdd FILL
XFILL_54_6 gnd vdd FILL
XFILL_3_INVX1_11 gnd vdd FILL
XFILL_63_2_2 gnd vdd FILL
XFILL_10_INVX8_1 gnd vdd FILL
XFILL_3_INVX1_22 gnd vdd FILL
XFILL_3_INVX1_33 gnd vdd FILL
XFILL_3_INVX1_44 gnd vdd FILL
XFILL_3_INVX1_55 gnd vdd FILL
XFILL_4_AND2X2_3 gnd vdd FILL
XFILL_3_INVX1_66 gnd vdd FILL
XFILL_3_INVX1_77 gnd vdd FILL
XFILL_49_DFFSR_14 gnd vdd FILL
XFILL_3_INVX1_88 gnd vdd FILL
XFILL_49_DFFSR_25 gnd vdd FILL
XFILL_3_INVX1_99 gnd vdd FILL
XFILL_49_DFFSR_36 gnd vdd FILL
XFILL_32_6_0 gnd vdd FILL
XFILL_49_DFFSR_47 gnd vdd FILL
XFILL_49_DFFSR_58 gnd vdd FILL
XFILL_49_DFFSR_69 gnd vdd FILL
XFILL_10_MUX2X1_9 gnd vdd FILL
XFILL_22_CLKBUF1_18 gnd vdd FILL
XFILL_1_BUFX4_20 gnd vdd FILL
XFILL_52_DFFSR_1 gnd vdd FILL
XFILL_1_BUFX4_31 gnd vdd FILL
XFILL_22_CLKBUF1_29 gnd vdd FILL
XFILL_1_BUFX4_42 gnd vdd FILL
XFILL_18_DFFSR_13 gnd vdd FILL
XFILL_18_DFFSR_24 gnd vdd FILL
XFILL_1_BUFX4_53 gnd vdd FILL
XFILL_1_BUFX4_64 gnd vdd FILL
XFILL_18_DFFSR_35 gnd vdd FILL
XFILL_1_BUFX4_75 gnd vdd FILL
XFILL_18_DFFSR_46 gnd vdd FILL
XFILL_1_BUFX4_86 gnd vdd FILL
XFILL_1_BUFX4_97 gnd vdd FILL
XFILL_13_DFFSR_101 gnd vdd FILL
XFILL_18_DFFSR_57 gnd vdd FILL
XFILL_18_DFFSR_68 gnd vdd FILL
XFILL_13_DFFSR_112 gnd vdd FILL
XFILL_18_DFFSR_79 gnd vdd FILL
XFILL_0_AOI21X1_19 gnd vdd FILL
XFILL_13_DFFSR_123 gnd vdd FILL
XFILL_13_DFFSR_134 gnd vdd FILL
XFILL_58_DFFSR_12 gnd vdd FILL
XFILL_13_DFFSR_145 gnd vdd FILL
XFILL_13_DFFSR_156 gnd vdd FILL
XFILL_58_DFFSR_23 gnd vdd FILL
XFILL_58_DFFSR_34 gnd vdd FILL
XFILL_29_NOR3X1_9 gnd vdd FILL
XFILL_13_DFFSR_167 gnd vdd FILL
XFILL_58_DFFSR_45 gnd vdd FILL
XFILL_13_DFFSR_178 gnd vdd FILL
XFILL_58_DFFSR_56 gnd vdd FILL
XFILL_17_DFFSR_100 gnd vdd FILL
XFILL_13_DFFSR_189 gnd vdd FILL
XFILL_58_DFFSR_67 gnd vdd FILL
XFILL_17_DFFSR_111 gnd vdd FILL
XFILL_58_DFFSR_78 gnd vdd FILL
XFILL_3_NOR2X1_107 gnd vdd FILL
XFILL_3_NOR2X1_118 gnd vdd FILL
XFILL_58_DFFSR_89 gnd vdd FILL
XFILL_17_DFFSR_122 gnd vdd FILL
XFILL_17_DFFSR_133 gnd vdd FILL
XFILL_4_DFFSR_6 gnd vdd FILL
XFILL_17_DFFSR_144 gnd vdd FILL
XFILL_3_NOR2X1_129 gnd vdd FILL
XFILL_17_DFFSR_155 gnd vdd FILL
XFILL_17_DFFSR_4 gnd vdd FILL
XFILL_17_DFFSR_166 gnd vdd FILL
XFILL_74_DFFSR_5 gnd vdd FILL
XFILL_6_CLKBUF1_9 gnd vdd FILL
XFILL_17_DFFSR_177 gnd vdd FILL
XFILL_27_DFFSR_11 gnd vdd FILL
XFILL_17_DFFSR_188 gnd vdd FILL
XFILL_27_DFFSR_22 gnd vdd FILL
XFILL_17_DFFSR_199 gnd vdd FILL
XFILL_27_DFFSR_33 gnd vdd FILL
XFILL_27_DFFSR_44 gnd vdd FILL
XFILL_27_DFFSR_55 gnd vdd FILL
XFILL_2_BUFX4_104 gnd vdd FILL
XFILL_27_DFFSR_66 gnd vdd FILL
XFILL_27_DFFSR_77 gnd vdd FILL
XFILL_27_DFFSR_88 gnd vdd FILL
XFILL_27_DFFSR_99 gnd vdd FILL
XFILL_13_NOR3X1_12 gnd vdd FILL
XFILL_67_DFFSR_10 gnd vdd FILL
XFILL_13_NOR3X1_23 gnd vdd FILL
XFILL_13_NOR3X1_34 gnd vdd FILL
XFILL_54_2_2 gnd vdd FILL
XFILL_67_DFFSR_21 gnd vdd FILL
XFILL_67_DFFSR_32 gnd vdd FILL
XFILL_63_DFFSR_201 gnd vdd FILL
XFILL_20_MUX2X1_109 gnd vdd FILL
XFILL_67_DFFSR_43 gnd vdd FILL
XFILL_2_MUX2X1_8 gnd vdd FILL
XFILL_13_NOR3X1_45 gnd vdd FILL
XFILL_63_DFFSR_212 gnd vdd FILL
XFILL_67_DFFSR_54 gnd vdd FILL
XFILL_67_DFFSR_65 gnd vdd FILL
XFILL_63_DFFSR_223 gnd vdd FILL
XFILL_63_DFFSR_234 gnd vdd FILL
XFILL_6_BUFX4_103 gnd vdd FILL
XFILL_67_DFFSR_76 gnd vdd FILL
XFILL_67_DFFSR_87 gnd vdd FILL
XFILL_63_DFFSR_245 gnd vdd FILL
XFILL_17_NOR3X1_11 gnd vdd FILL
XFILL_67_DFFSR_98 gnd vdd FILL
XFILL_63_DFFSR_256 gnd vdd FILL
XFILL_63_DFFSR_267 gnd vdd FILL
XFILL_23_6_0 gnd vdd FILL
XFILL_17_NOR3X1_22 gnd vdd FILL
XFILL_17_NOR3X1_33 gnd vdd FILL
XFILL_17_NOR3X1_44 gnd vdd FILL
XFILL_67_DFFSR_200 gnd vdd FILL
XFILL_67_DFFSR_211 gnd vdd FILL
XFILL_39_DFFSR_8 gnd vdd FILL
XFILL_67_DFFSR_222 gnd vdd FILL
XFILL_36_DFFSR_20 gnd vdd FILL
XFILL_67_DFFSR_233 gnd vdd FILL
XFILL_0_OAI22X1_16 gnd vdd FILL
XFILL_36_DFFSR_31 gnd vdd FILL
XFILL_0_OAI22X1_27 gnd vdd FILL
XFILL_36_DFFSR_42 gnd vdd FILL
XFILL_67_DFFSR_244 gnd vdd FILL
XFILL_67_DFFSR_255 gnd vdd FILL
XFILL_36_DFFSR_53 gnd vdd FILL
XFILL_0_OAI22X1_38 gnd vdd FILL
XFILL_36_DFFSR_64 gnd vdd FILL
XFILL_67_DFFSR_266 gnd vdd FILL
XFILL_0_OAI22X1_49 gnd vdd FILL
XFILL_22_CLKBUF1_7 gnd vdd FILL
XFILL_36_DFFSR_75 gnd vdd FILL
XAOI21X1_10 BUFX4_74/Y AOI21X1_9/B NOR2X1_146/Y gnd DFFSR_105/D vdd AOI21X1
XFILL_4_OAI21X1_18 gnd vdd FILL
XAOI21X1_21 MUX2X1_66/A MUX2X1_9/S NOR2X1_173/Y gnd DFFSR_40/D vdd AOI21X1
XFILL_4_OAI21X1_29 gnd vdd FILL
XFILL_36_DFFSR_86 gnd vdd FILL
XFILL_36_DFFSR_97 gnd vdd FILL
XFILL_0_NOR2X1_17 gnd vdd FILL
XAOI21X1_32 BUFX4_78/Y NOR2X1_190/B NOR2X1_189/Y gnd DFFSR_21/D vdd AOI21X1
XFILL_0_NOR2X1_28 gnd vdd FILL
XAOI21X1_43 BUFX4_85/Y MUX2X1_22/S NOR2X1_204/Y gnd DFFSR_275/D vdd AOI21X1
XFILL_76_DFFSR_30 gnd vdd FILL
XFILL_0_NOR2X1_39 gnd vdd FILL
XAOI21X1_54 BUFX4_85/Y NOR2X1_16/B NOR2X1_15/Y gnd DFFSR_258/D vdd AOI21X1
XFILL_76_DFFSR_41 gnd vdd FILL
XAOI21X1_65 NAND3X1_67/Y OAI21X1_23/Y NOR3X1_9/A gnd AND2X2_6/A vdd AOI21X1
XAOI21X1_76 OAI21X1_41/A INVX1_57/A AOI22X1_3/A gnd NOR3X1_48/C vdd AOI21X1
XFILL_76_DFFSR_52 gnd vdd FILL
XFILL_76_DFFSR_63 gnd vdd FILL
XFILL_76_DFFSR_74 gnd vdd FILL
XFILL_26_CLKBUF1_6 gnd vdd FILL
XFILL_76_DFFSR_85 gnd vdd FILL
XFILL_3_NAND2X1_50 gnd vdd FILL
XFILL_4_NOR2X1_16 gnd vdd FILL
XOAI21X1_5 OAI21X1_5/A OAI21X1_5/B OAI21X1_5/C gnd OAI21X1_5/Y vdd OAI21X1
XFILL_76_DFFSR_96 gnd vdd FILL
XFILL_3_NAND2X1_61 gnd vdd FILL
XFILL_11_BUFX4_4 gnd vdd FILL
XFILL_4_NOR2X1_27 gnd vdd FILL
XFILL_3_NAND2X1_72 gnd vdd FILL
XFILL_3_NAND2X1_83 gnd vdd FILL
XFILL_4_NOR2X1_38 gnd vdd FILL
XFILL_4_NOR2X1_49 gnd vdd FILL
XFILL_3_NAND2X1_94 gnd vdd FILL
XFILL_45_DFFSR_40 gnd vdd FILL
XFILL_11_CLKBUF1_14 gnd vdd FILL
XFILL_16_NOR3X1_4 gnd vdd FILL
XFILL_8_NOR2X1_15 gnd vdd FILL
XFILL_8_NOR2X1_26 gnd vdd FILL
XFILL_11_CLKBUF1_25 gnd vdd FILL
XFILL_45_DFFSR_51 gnd vdd FILL
XFILL_11_CLKBUF1_36 gnd vdd FILL
XFILL_45_DFFSR_62 gnd vdd FILL
XFILL_8_NOR2X1_37 gnd vdd FILL
XFILL_45_DFFSR_73 gnd vdd FILL
XFILL_6_7_0 gnd vdd FILL
XFILL_45_DFFSR_84 gnd vdd FILL
XFILL_8_NOR2X1_48 gnd vdd FILL
XFILL_45_DFFSR_95 gnd vdd FILL
XFILL_8_NOR2X1_59 gnd vdd FILL
XFILL_85_DFFSR_50 gnd vdd FILL
XFILL_85_DFFSR_61 gnd vdd FILL
XFILL_85_DFFSR_72 gnd vdd FILL
XFILL_85_DFFSR_83 gnd vdd FILL
XFILL_45_2_2 gnd vdd FILL
XFILL_85_DFFSR_94 gnd vdd FILL
XFILL_16_OAI22X1_9 gnd vdd FILL
XFILL_14_DFFSR_50 gnd vdd FILL
XFILL_14_DFFSR_61 gnd vdd FILL
XFILL_14_DFFSR_72 gnd vdd FILL
XFILL_14_DFFSR_83 gnd vdd FILL
XFILL_14_DFFSR_94 gnd vdd FILL
XFILL_30_DFFSR_201 gnd vdd FILL
XFILL_30_DFFSR_212 gnd vdd FILL
XFILL_30_DFFSR_223 gnd vdd FILL
XFILL_14_6_0 gnd vdd FILL
XFILL_25_NOR3X1_2 gnd vdd FILL
XFILL_30_DFFSR_234 gnd vdd FILL
XFILL_30_DFFSR_245 gnd vdd FILL
XFILL_54_DFFSR_60 gnd vdd FILL
XOAI22X1_40 INVX1_187/Y OAI22X1_50/B INVX1_182/Y OAI22X1_50/D gnd OAI22X1_40/Y vdd
+ OAI22X1
XOAI22X1_51 MUX2X1_92/A OAI22X1_7/D MUX2X1_96/A NOR2X1_60/B gnd OAI22X1_51/Y vdd OAI22X1
XFILL_7_AOI21X1_50 gnd vdd FILL
XFILL_30_DFFSR_256 gnd vdd FILL
XFILL_30_DFFSR_267 gnd vdd FILL
XFILL_54_DFFSR_71 gnd vdd FILL
XFILL_7_AOI21X1_61 gnd vdd FILL
XFILL_54_DFFSR_82 gnd vdd FILL
XFILL_7_AOI21X1_72 gnd vdd FILL
XFILL_54_DFFSR_93 gnd vdd FILL
XFILL_17_OAI22X1_30 gnd vdd FILL
XFILL_17_OAI22X1_41 gnd vdd FILL
XFILL_34_DFFSR_200 gnd vdd FILL
XFILL_34_DFFSR_211 gnd vdd FILL
XFILL_34_DFFSR_222 gnd vdd FILL
XFILL_34_DFFSR_233 gnd vdd FILL
XFILL_34_DFFSR_244 gnd vdd FILL
XFILL_34_DFFSR_255 gnd vdd FILL
XFILL_1_CLKBUF1_20 gnd vdd FILL
XFILL_0_MUX2X1_13 gnd vdd FILL
XFILL_34_DFFSR_266 gnd vdd FILL
XFILL_1_CLKBUF1_31 gnd vdd FILL
XFILL_61_DFFSR_100 gnd vdd FILL
XFILL_1_CLKBUF1_42 gnd vdd FILL
XFILL_0_MUX2X1_24 gnd vdd FILL
XFILL_1_INVX8_4 gnd vdd FILL
XFILL_0_MUX2X1_35 gnd vdd FILL
XFILL_61_DFFSR_111 gnd vdd FILL
XFILL_38_DFFSR_210 gnd vdd FILL
XFILL_23_DFFSR_70 gnd vdd FILL
XFILL_0_MUX2X1_46 gnd vdd FILL
XFILL_14_INVX8_2 gnd vdd FILL
XFILL_38_DFFSR_221 gnd vdd FILL
XFILL_0_MUX2X1_57 gnd vdd FILL
XFILL_61_DFFSR_122 gnd vdd FILL
XFILL_61_DFFSR_133 gnd vdd FILL
XFILL_0_MUX2X1_68 gnd vdd FILL
XFILL_38_DFFSR_232 gnd vdd FILL
XFILL_23_DFFSR_81 gnd vdd FILL
XFILL_38_DFFSR_243 gnd vdd FILL
XFILL_23_DFFSR_92 gnd vdd FILL
XFILL_61_DFFSR_144 gnd vdd FILL
XFILL_0_MUX2X1_79 gnd vdd FILL
XFILL_61_DFFSR_155 gnd vdd FILL
XFILL_8_NOR3X1_3 gnd vdd FILL
XFILL_38_DFFSR_254 gnd vdd FILL
XFILL_61_DFFSR_166 gnd vdd FILL
XFILL_4_MUX2X1_12 gnd vdd FILL
XFILL_38_DFFSR_265 gnd vdd FILL
XFILL_4_MUX2X1_23 gnd vdd FILL
XFILL_61_DFFSR_177 gnd vdd FILL
XFILL_61_DFFSR_188 gnd vdd FILL
XFILL_4_MUX2X1_34 gnd vdd FILL
XFILL_65_DFFSR_110 gnd vdd FILL
XFILL_61_DFFSR_199 gnd vdd FILL
XFILL_10_OAI21X1_10 gnd vdd FILL
XFILL_4_MUX2X1_45 gnd vdd FILL
XFILL_65_DFFSR_121 gnd vdd FILL
XFILL_63_DFFSR_80 gnd vdd FILL
XFILL_10_OAI21X1_21 gnd vdd FILL
XFILL_4_MUX2X1_56 gnd vdd FILL
XFILL_65_DFFSR_132 gnd vdd FILL
XFILL_10_OAI21X1_32 gnd vdd FILL
XFILL_4_MUX2X1_67 gnd vdd FILL
XFILL_65_DFFSR_143 gnd vdd FILL
XFILL_63_DFFSR_91 gnd vdd FILL
XFILL_10_OAI21X1_43 gnd vdd FILL
XFILL_65_DFFSR_154 gnd vdd FILL
XFILL_4_MUX2X1_78 gnd vdd FILL
XFILL_3_2 gnd vdd FILL
XFILL_65_DFFSR_165 gnd vdd FILL
XFILL_4_MUX2X1_89 gnd vdd FILL
XFILL_8_MUX2X1_11 gnd vdd FILL
XFILL_8_MUX2X1_22 gnd vdd FILL
XFILL_65_DFFSR_176 gnd vdd FILL
XFILL_65_DFFSR_187 gnd vdd FILL
XFILL_8_MUX2X1_33 gnd vdd FILL
XFILL_65_DFFSR_198 gnd vdd FILL
XFILL_56_DFFSR_2 gnd vdd FILL
XFILL_69_DFFSR_120 gnd vdd FILL
XFILL_8_MUX2X1_44 gnd vdd FILL
XFILL_69_DFFSR_131 gnd vdd FILL
XFILL_8_MUX2X1_55 gnd vdd FILL
XFILL_6_DFFSR_60 gnd vdd FILL
XFILL_8_MUX2X1_66 gnd vdd FILL
XFILL_6_DFFSR_71 gnd vdd FILL
XFILL_8_MUX2X1_77 gnd vdd FILL
XFILL_69_DFFSR_142 gnd vdd FILL
XFILL_6_DFFSR_82 gnd vdd FILL
XFILL_69_DFFSR_153 gnd vdd FILL
XFILL_8_MUX2X1_88 gnd vdd FILL
XFILL_6_DFFSR_93 gnd vdd FILL
XFILL_69_DFFSR_164 gnd vdd FILL
XFILL_8_MUX2X1_99 gnd vdd FILL
XFILL_69_DFFSR_175 gnd vdd FILL
XFILL_64_5_0 gnd vdd FILL
XFILL_32_DFFSR_90 gnd vdd FILL
XFILL_69_DFFSR_186 gnd vdd FILL
XFILL_36_2_2 gnd vdd FILL
XFILL_69_DFFSR_197 gnd vdd FILL
XFILL_45_2 gnd vdd FILL
XFILL_38_1 gnd vdd FILL
XFILL_20_MUX2X1_10 gnd vdd FILL
XFILL_20_MUX2X1_21 gnd vdd FILL
XFILL_40_DFFSR_8 gnd vdd FILL
XFILL_20_MUX2X1_32 gnd vdd FILL
XFILL_8_DFFSR_7 gnd vdd FILL
XFILL_20_MUX2X1_43 gnd vdd FILL
XFILL_20_MUX2X1_54 gnd vdd FILL
XFILL_12_NAND3X1_19 gnd vdd FILL
XFILL_20_MUX2X1_65 gnd vdd FILL
XFILL_20_MUX2X1_76 gnd vdd FILL
XFILL_78_DFFSR_6 gnd vdd FILL
XFILL_20_MUX2X1_87 gnd vdd FILL
XFILL_20_MUX2X1_98 gnd vdd FILL
XFILL_32_CLKBUF1_19 gnd vdd FILL
XFILL_32_DFFSR_110 gnd vdd FILL
XFILL_32_DFFSR_121 gnd vdd FILL
XFILL_32_DFFSR_132 gnd vdd FILL
XFILL_32_DFFSR_143 gnd vdd FILL
XFILL_32_DFFSR_154 gnd vdd FILL
XFILL_32_DFFSR_165 gnd vdd FILL
XFILL_32_DFFSR_176 gnd vdd FILL
XFILL_32_DFFSR_187 gnd vdd FILL
XFILL_32_DFFSR_198 gnd vdd FILL
XFILL_36_DFFSR_120 gnd vdd FILL
XFILL_2_NAND3X1_14 gnd vdd FILL
XFILL_36_DFFSR_131 gnd vdd FILL
XFILL_2_NAND3X1_25 gnd vdd FILL
XFILL_55_5_0 gnd vdd FILL
XFILL_36_DFFSR_142 gnd vdd FILL
XFILL_2_NAND3X1_36 gnd vdd FILL
XFILL_36_DFFSR_153 gnd vdd FILL
XFILL_2_NAND3X1_47 gnd vdd FILL
XFILL_27_2_2 gnd vdd FILL
XFILL_2_NAND3X1_58 gnd vdd FILL
XFILL_2_2_2 gnd vdd FILL
XFILL_36_DFFSR_164 gnd vdd FILL
XFILL_36_DFFSR_175 gnd vdd FILL
XFILL_6_NAND2X1_16 gnd vdd FILL
XFILL_2_NAND3X1_69 gnd vdd FILL
XFILL_6_NAND2X1_27 gnd vdd FILL
XFILL_36_DFFSR_186 gnd vdd FILL
XFILL_6_NAND2X1_38 gnd vdd FILL
XFILL_36_DFFSR_197 gnd vdd FILL
XFILL_2_BUFX4_7 gnd vdd FILL
XFILL_6_NAND2X1_49 gnd vdd FILL
XFILL_15_BUFX4_5 gnd vdd FILL
XMUX2X1_9 MUX2X1_9/A MUX2X1_9/B MUX2X1_9/S gnd MUX2X1_9/Y vdd MUX2X1
XFILL_16_MUX2X1_180 gnd vdd FILL
XFILL_16_MUX2X1_191 gnd vdd FILL
XFILL_82_DFFSR_210 gnd vdd FILL
XFILL_82_DFFSR_221 gnd vdd FILL
XFILL_82_DFFSR_232 gnd vdd FILL
XFILL_10_1_2 gnd vdd FILL
XFILL_82_DFFSR_243 gnd vdd FILL
XFILL_82_DFFSR_254 gnd vdd FILL
XFILL_82_DFFSR_265 gnd vdd FILL
XFILL_18_DFFSR_109 gnd vdd FILL
XFILL_86_DFFSR_220 gnd vdd FILL
XFILL_13_AOI21X1_5 gnd vdd FILL
XFILL_86_DFFSR_231 gnd vdd FILL
XFILL_86_DFFSR_242 gnd vdd FILL
XFILL_86_DFFSR_253 gnd vdd FILL
XFILL_86_DFFSR_264 gnd vdd FILL
XFILL_86_DFFSR_275 gnd vdd FILL
XFILL_11_BUFX2_1 gnd vdd FILL
XFILL_2_INVX1_170 gnd vdd FILL
XFILL_2_INVX1_181 gnd vdd FILL
XFILL_77_DFFSR_19 gnd vdd FILL
XFILL_2_INVX1_192 gnd vdd FILL
XFILL_21_CLKBUF1_15 gnd vdd FILL
XFILL_21_CLKBUF1_26 gnd vdd FILL
XBUFX4_104 BUFX4_2/A gnd BUFX4_104/Y vdd BUFX4
XFILL_21_CLKBUF1_37 gnd vdd FILL
XFILL_0_INVX1_15 gnd vdd FILL
XFILL_6_INVX1_180 gnd vdd FILL
XFILL_0_INVX1_26 gnd vdd FILL
XFILL_4_CLKBUF1_19 gnd vdd FILL
XFILL_0_INVX1_37 gnd vdd FILL
XFILL_6_INVX1_191 gnd vdd FILL
XFILL_46_5_0 gnd vdd FILL
XFILL_0_INVX1_48 gnd vdd FILL
XFILL_1_AND2X2_7 gnd vdd FILL
XFILL_18_2_2 gnd vdd FILL
XFILL_0_INVX1_59 gnd vdd FILL
XFILL_68_DFFSR_209 gnd vdd FILL
XFILL_18_INVX8_3 gnd vdd FILL
XFILL_46_DFFSR_18 gnd vdd FILL
XFILL_46_DFFSR_29 gnd vdd FILL
XFILL_31_8 gnd vdd FILL
XFILL_60_0_2 gnd vdd FILL
XFILL_2_NOR2X1_104 gnd vdd FILL
XFILL_24_7 gnd vdd FILL
XFILL_2_NOR2X1_115 gnd vdd FILL
XFILL_2_NOR2X1_126 gnd vdd FILL
XFILL_86_DFFSR_17 gnd vdd FILL
XFILL_86_DFFSR_28 gnd vdd FILL
XFILL_22_DFFSR_5 gnd vdd FILL
XFILL_86_DFFSR_39 gnd vdd FILL
XFILL_2_NOR2X1_137 gnd vdd FILL
XFILL_2_NOR2X1_148 gnd vdd FILL
XFILL_2_NOR2X1_159 gnd vdd FILL
XFILL_15_DFFSR_17 gnd vdd FILL
XFILL_15_DFFSR_28 gnd vdd FILL
XFILL_15_DFFSR_39 gnd vdd FILL
XFILL_55_DFFSR_16 gnd vdd FILL
XFILL_55_DFFSR_27 gnd vdd FILL
XFILL_55_DFFSR_38 gnd vdd FILL
XFILL_55_DFFSR_49 gnd vdd FILL
XFILL_53_DFFSR_220 gnd vdd FILL
XFILL_53_DFFSR_231 gnd vdd FILL
XFILL_53_DFFSR_242 gnd vdd FILL
XFILL_53_DFFSR_253 gnd vdd FILL
XFILL_53_DFFSR_264 gnd vdd FILL
XFILL_53_DFFSR_275 gnd vdd FILL
XFILL_44_DFFSR_9 gnd vdd FILL
XFILL_80_DFFSR_120 gnd vdd FILL
XFILL_24_DFFSR_15 gnd vdd FILL
XFILL_7_NOR2X1_204 gnd vdd FILL
XFILL_24_DFFSR_26 gnd vdd FILL
XFILL_80_DFFSR_131 gnd vdd FILL
XFILL_24_DFFSR_37 gnd vdd FILL
XFILL_57_DFFSR_230 gnd vdd FILL
XFILL_80_DFFSR_142 gnd vdd FILL
XFILL_57_DFFSR_241 gnd vdd FILL
XFILL_24_DFFSR_48 gnd vdd FILL
XFILL_15_BUFX4_80 gnd vdd FILL
XFILL_80_DFFSR_153 gnd vdd FILL
XFILL_24_DFFSR_59 gnd vdd FILL
XFILL_15_BUFX4_91 gnd vdd FILL
XFILL_57_DFFSR_252 gnd vdd FILL
XFILL_80_DFFSR_164 gnd vdd FILL
XFILL_57_DFFSR_263 gnd vdd FILL
XFILL_57_DFFSR_274 gnd vdd FILL
XFILL_3_OAI21X1_15 gnd vdd FILL
XFILL_80_DFFSR_175 gnd vdd FILL
XFILL_12_CLKBUF1_4 gnd vdd FILL
XFILL_0_DFFSR_201 gnd vdd FILL
XFILL_80_DFFSR_186 gnd vdd FILL
XFILL_3_OAI21X1_26 gnd vdd FILL
XFILL_80_DFFSR_197 gnd vdd FILL
XFILL_0_DFFSR_212 gnd vdd FILL
XFILL_64_DFFSR_14 gnd vdd FILL
XFILL_0_DFFSR_223 gnd vdd FILL
XFILL_3_OAI21X1_37 gnd vdd FILL
XFILL_0_DFFSR_234 gnd vdd FILL
XFILL_64_DFFSR_25 gnd vdd FILL
XFILL_3_OAI21X1_48 gnd vdd FILL
XFILL_84_DFFSR_130 gnd vdd FILL
XFILL_64_DFFSR_36 gnd vdd FILL
XFILL_37_5_0 gnd vdd FILL
XFILL_0_DFFSR_245 gnd vdd FILL
XFILL_84_DFFSR_141 gnd vdd FILL
XFILL_64_DFFSR_47 gnd vdd FILL
XFILL_84_DFFSR_152 gnd vdd FILL
XFILL_64_DFFSR_58 gnd vdd FILL
XFILL_0_DFFSR_256 gnd vdd FILL
XFILL_0_DFFSR_267 gnd vdd FILL
XFILL_64_DFFSR_69 gnd vdd FILL
XFILL_84_DFFSR_163 gnd vdd FILL
XFILL_84_DFFSR_174 gnd vdd FILL
XFILL_16_CLKBUF1_3 gnd vdd FILL
XFILL_4_DFFSR_200 gnd vdd FILL
XFILL_84_DFFSR_185 gnd vdd FILL
XFILL_4_DFFSR_211 gnd vdd FILL
XFILL_84_DFFSR_196 gnd vdd FILL
XFILL_4_DFFSR_222 gnd vdd FILL
XFILL_35_DFFSR_209 gnd vdd FILL
XFILL_4_DFFSR_233 gnd vdd FILL
XFILL_2_NAND2X1_80 gnd vdd FILL
XFILL_7_DFFSR_16 gnd vdd FILL
XFILL_2_NAND2X1_91 gnd vdd FILL
XFILL_7_DFFSR_27 gnd vdd FILL
XFILL_4_DFFSR_244 gnd vdd FILL
XFILL_33_DFFSR_13 gnd vdd FILL
XFILL_51_0_2 gnd vdd FILL
XFILL_4_DFFSR_255 gnd vdd FILL
XFILL_7_DFFSR_38 gnd vdd FILL
XFILL_33_DFFSR_24 gnd vdd FILL
XFILL_7_DFFSR_49 gnd vdd FILL
XFILL_4_DFFSR_266 gnd vdd FILL
XFILL_33_DFFSR_35 gnd vdd FILL
XFILL_10_CLKBUF1_11 gnd vdd FILL
XFILL_33_DFFSR_46 gnd vdd FILL
XFILL_10_CLKBUF1_22 gnd vdd FILL
XFILL_62_DFFSR_109 gnd vdd FILL
XFILL_8_DFFSR_210 gnd vdd FILL
XFILL_33_DFFSR_57 gnd vdd FILL
XFILL_39_DFFSR_208 gnd vdd FILL
XFILL_33_DFFSR_68 gnd vdd FILL
XFILL_8_DFFSR_221 gnd vdd FILL
XFILL_39_DFFSR_219 gnd vdd FILL
XFILL_10_CLKBUF1_33 gnd vdd FILL
XFILL_33_DFFSR_79 gnd vdd FILL
XFILL_8_DFFSR_232 gnd vdd FILL
XFILL_8_DFFSR_243 gnd vdd FILL
XFILL_20_4_0 gnd vdd FILL
XFILL_73_DFFSR_12 gnd vdd FILL
XFILL_8_DFFSR_254 gnd vdd FILL
XFILL_73_DFFSR_23 gnd vdd FILL
XFILL_8_DFFSR_265 gnd vdd FILL
XFILL_73_DFFSR_34 gnd vdd FILL
XFILL_16_MUX2X1_2 gnd vdd FILL
XFILL_73_DFFSR_45 gnd vdd FILL
XFILL_73_DFFSR_56 gnd vdd FILL
XFILL_66_DFFSR_108 gnd vdd FILL
XFILL_73_DFFSR_67 gnd vdd FILL
XFILL_66_DFFSR_119 gnd vdd FILL
XFILL_73_DFFSR_78 gnd vdd FILL
XFILL_73_DFFSR_89 gnd vdd FILL
XFILL_6_BUFX4_8 gnd vdd FILL
XFILL_42_DFFSR_11 gnd vdd FILL
XFILL_42_DFFSR_22 gnd vdd FILL
XFILL_19_MUX2X1_102 gnd vdd FILL
XFILL_10_NOR2X1_11 gnd vdd FILL
XFILL_42_DFFSR_33 gnd vdd FILL
XFILL_13_NOR3X1_8 gnd vdd FILL
XFILL_19_MUX2X1_113 gnd vdd FILL
XFILL_7_BUFX4_90 gnd vdd FILL
XFILL_20_DFFSR_220 gnd vdd FILL
XFILL_10_NOR2X1_22 gnd vdd FILL
XFILL_42_DFFSR_44 gnd vdd FILL
XFILL_19_MUX2X1_124 gnd vdd FILL
XFILL_1_AOI22X1_5 gnd vdd FILL
XFILL_20_DFFSR_231 gnd vdd FILL
XFILL_42_DFFSR_55 gnd vdd FILL
XFILL_13_OAI21X1_8 gnd vdd FILL
XFILL_10_NOR2X1_33 gnd vdd FILL
XFILL_20_DFFSR_242 gnd vdd FILL
XFILL_10_NOR2X1_44 gnd vdd FILL
XFILL_19_MUX2X1_135 gnd vdd FILL
XFILL_42_DFFSR_66 gnd vdd FILL
XFILL_42_DFFSR_77 gnd vdd FILL
XFILL_10_NOR2X1_55 gnd vdd FILL
XFILL_19_MUX2X1_146 gnd vdd FILL
XFILL_20_DFFSR_253 gnd vdd FILL
XFILL_10_NOR2X1_66 gnd vdd FILL
XFILL_42_DFFSR_88 gnd vdd FILL
XFILL_20_DFFSR_264 gnd vdd FILL
XFILL_19_MUX2X1_157 gnd vdd FILL
XFILL_20_DFFSR_275 gnd vdd FILL
XFILL_42_DFFSR_99 gnd vdd FILL
XFILL_19_MUX2X1_168 gnd vdd FILL
XFILL_10_NOR2X1_77 gnd vdd FILL
XFILL_1_INVX1_204 gnd vdd FILL
XFILL_6_AOI21X1_80 gnd vdd FILL
XFILL_82_DFFSR_10 gnd vdd FILL
XFILL_19_MUX2X1_179 gnd vdd FILL
XFILL_59_1_2 gnd vdd FILL
XFILL_82_DFFSR_21 gnd vdd FILL
XFILL_1_INVX1_215 gnd vdd FILL
XFILL_10_NOR2X1_88 gnd vdd FILL
XFILL_10_NOR2X1_99 gnd vdd FILL
XFILL_82_DFFSR_32 gnd vdd FILL
XFILL_1_INVX1_226 gnd vdd FILL
XFILL_82_DFFSR_43 gnd vdd FILL
XFILL_24_DFFSR_230 gnd vdd FILL
XFILL_11_DFFSR_10 gnd vdd FILL
XFILL_82_DFFSR_54 gnd vdd FILL
XFILL_5_AOI22X1_4 gnd vdd FILL
XFILL_24_DFFSR_241 gnd vdd FILL
XFILL_11_DFFSR_21 gnd vdd FILL
XFILL_82_DFFSR_65 gnd vdd FILL
XFILL_82_DFFSR_76 gnd vdd FILL
XFILL_24_DFFSR_252 gnd vdd FILL
XFILL_11_DFFSR_32 gnd vdd FILL
XFILL_11_DFFSR_43 gnd vdd FILL
XFILL_82_DFFSR_87 gnd vdd FILL
XFILL_24_DFFSR_263 gnd vdd FILL
XFILL_24_DFFSR_274 gnd vdd FILL
XFILL_82_DFFSR_98 gnd vdd FILL
XFILL_11_DFFSR_54 gnd vdd FILL
XFILL_28_5_0 gnd vdd FILL
XFILL_21_MUX2X1_19 gnd vdd FILL
XFILL_5_INVX1_203 gnd vdd FILL
XFILL_3_5_0 gnd vdd FILL
XFILL_9_NOR2X1_3 gnd vdd FILL
XFILL_11_DFFSR_65 gnd vdd FILL
XFILL_9_NOR2X1_190 gnd vdd FILL
XFILL_5_INVX1_214 gnd vdd FILL
XFILL_11_DFFSR_76 gnd vdd FILL
XFILL_5_INVX1_225 gnd vdd FILL
XFILL_11_DFFSR_87 gnd vdd FILL
XFILL_51_DFFSR_130 gnd vdd FILL
XFILL_11_DFFSR_98 gnd vdd FILL
XFILL_9_AOI22X1_3 gnd vdd FILL
XFILL_28_DFFSR_240 gnd vdd FILL
XFILL_51_DFFSR_141 gnd vdd FILL
XFILL_51_DFFSR_152 gnd vdd FILL
XFILL_28_DFFSR_251 gnd vdd FILL
XFILL_51_DFFSR_20 gnd vdd FILL
XFILL_51_DFFSR_163 gnd vdd FILL
XFILL_51_DFFSR_31 gnd vdd FILL
XFILL_51_DFFSR_174 gnd vdd FILL
XFILL_2_BUFX2_4 gnd vdd FILL
XFILL_22_NOR3X1_6 gnd vdd FILL
XFILL_28_DFFSR_262 gnd vdd FILL
XFILL_51_DFFSR_42 gnd vdd FILL
XFILL_51_DFFSR_53 gnd vdd FILL
XFILL_28_DFFSR_273 gnd vdd FILL
XFILL_51_DFFSR_64 gnd vdd FILL
XFILL_51_DFFSR_185 gnd vdd FILL
XFILL_42_0_2 gnd vdd FILL
XFILL_51_DFFSR_196 gnd vdd FILL
XFILL_51_DFFSR_75 gnd vdd FILL
XFILL_51_DFFSR_86 gnd vdd FILL
XFILL_51_DFFSR_97 gnd vdd FILL
XFILL_55_DFFSR_140 gnd vdd FILL
XFILL_8_MUX2X1_1 gnd vdd FILL
XFILL_55_DFFSR_151 gnd vdd FILL
XFILL_55_DFFSR_162 gnd vdd FILL
XFILL_55_DFFSR_173 gnd vdd FILL
XFILL_55_DFFSR_184 gnd vdd FILL
XFILL_11_4_0 gnd vdd FILL
XFILL_61_DFFSR_3 gnd vdd FILL
XFILL_55_DFFSR_195 gnd vdd FILL
XFILL_20_DFFSR_30 gnd vdd FILL
XFILL_20_DFFSR_41 gnd vdd FILL
XFILL_9_MUX2X1_130 gnd vdd FILL
XFILL_9_MUX2X1_141 gnd vdd FILL
XFILL_20_DFFSR_52 gnd vdd FILL
XFILL_20_DFFSR_63 gnd vdd FILL
XFILL_9_MUX2X1_152 gnd vdd FILL
XFILL_59_DFFSR_150 gnd vdd FILL
XFILL_20_DFFSR_74 gnd vdd FILL
XFILL_59_DFFSR_161 gnd vdd FILL
XFILL_9_MUX2X1_163 gnd vdd FILL
XFILL_59_DFFSR_172 gnd vdd FILL
XFILL_20_DFFSR_85 gnd vdd FILL
XFILL_9_MUX2X1_174 gnd vdd FILL
XFILL_9_MUX2X1_185 gnd vdd FILL
XFILL_59_DFFSR_183 gnd vdd FILL
XFILL_20_DFFSR_96 gnd vdd FILL
XFILL_2_DFFSR_110 gnd vdd FILL
XFILL_5_NOR3X1_7 gnd vdd FILL
XFILL_33_DFFSR_108 gnd vdd FILL
XFILL_59_DFFSR_194 gnd vdd FILL
XFILL_2_DFFSR_121 gnd vdd FILL
XFILL_33_DFFSR_119 gnd vdd FILL
XFILL_31_NOR3X1_4 gnd vdd FILL
XFILL_60_DFFSR_40 gnd vdd FILL
XFILL_2_DFFSR_132 gnd vdd FILL
XFILL_60_DFFSR_51 gnd vdd FILL
XFILL_2_DFFSR_143 gnd vdd FILL
XFILL_2_DFFSR_154 gnd vdd FILL
XFILL_60_DFFSR_62 gnd vdd FILL
XFILL_2_DFFSR_165 gnd vdd FILL
XFILL_60_DFFSR_73 gnd vdd FILL
XFILL_60_DFFSR_84 gnd vdd FILL
XFILL_2_DFFSR_176 gnd vdd FILL
XFILL_60_DFFSR_95 gnd vdd FILL
XFILL_2_DFFSR_187 gnd vdd FILL
XFILL_2_DFFSR_198 gnd vdd FILL
XFILL_37_DFFSR_107 gnd vdd FILL
XFILL_6_DFFSR_120 gnd vdd FILL
XFILL_6_DFFSR_131 gnd vdd FILL
XFILL_3_DFFSR_20 gnd vdd FILL
XFILL_37_DFFSR_118 gnd vdd FILL
XFILL_6_DFFSR_142 gnd vdd FILL
XFILL_10_MUX2X1_40 gnd vdd FILL
XFILL_3_DFFSR_31 gnd vdd FILL
XFILL_37_DFFSR_129 gnd vdd FILL
XFILL_6_DFFSR_153 gnd vdd FILL
XFILL_10_MUX2X1_51 gnd vdd FILL
XFILL_26_DFFSR_6 gnd vdd FILL
XFILL_3_DFFSR_42 gnd vdd FILL
XFILL_11_NAND3X1_16 gnd vdd FILL
XFILL_10_MUX2X1_62 gnd vdd FILL
XFILL_3_DFFSR_53 gnd vdd FILL
XFILL_6_DFFSR_164 gnd vdd FILL
XFILL_10_MUX2X1_73 gnd vdd FILL
XFILL_6_DFFSR_175 gnd vdd FILL
XFILL_11_NAND3X1_27 gnd vdd FILL
XFILL_3_DFFSR_64 gnd vdd FILL
XFILL_83_DFFSR_7 gnd vdd FILL
XFILL_3_DFFSR_75 gnd vdd FILL
XFILL_11_NAND3X1_38 gnd vdd FILL
XFILL_10_MUX2X1_84 gnd vdd FILL
XFILL_6_DFFSR_186 gnd vdd FILL
XFILL_6_DFFSR_197 gnd vdd FILL
XFILL_3_DFFSR_86 gnd vdd FILL
XFILL_10_MUX2X1_95 gnd vdd FILL
XFILL_11_NAND3X1_49 gnd vdd FILL
XFILL_2_INVX2_4 gnd vdd FILL
XFILL_3_DFFSR_97 gnd vdd FILL
XFILL_31_CLKBUF1_16 gnd vdd FILL
XFILL_31_CLKBUF1_27 gnd vdd FILL
XFILL_31_CLKBUF1_38 gnd vdd FILL
XFILL_14_MUX2X1_50 gnd vdd FILL
XFILL_14_MUX2X1_61 gnd vdd FILL
XFILL_19_5_0 gnd vdd FILL
XFILL_14_MUX2X1_72 gnd vdd FILL
XFILL_2_NOR3X1_10 gnd vdd FILL
XFILL_14_MUX2X1_83 gnd vdd FILL
XFILL_2_NOR3X1_21 gnd vdd FILL
XFILL_14_MUX2X1_94 gnd vdd FILL
XFILL_2_NOR3X1_32 gnd vdd FILL
XFILL_2_NOR3X1_43 gnd vdd FILL
XFILL_83_DFFSR_208 gnd vdd FILL
XFILL_83_DFFSR_219 gnd vdd FILL
XFILL_61_3_0 gnd vdd FILL
XFILL_0_INVX1_2 gnd vdd FILL
XFILL_18_MUX2X1_60 gnd vdd FILL
XFILL_18_MUX2X1_71 gnd vdd FILL
XFILL_33_0_2 gnd vdd FILL
XFILL_18_MUX2X1_82 gnd vdd FILL
XFILL_22_4 gnd vdd FILL
XFILL_6_NOR3X1_20 gnd vdd FILL
XFILL_18_MUX2X1_93 gnd vdd FILL
XFILL_6_NOR3X1_31 gnd vdd FILL
XFILL_6_NOR3X1_42 gnd vdd FILL
XFILL_87_DFFSR_207 gnd vdd FILL
XFILL_15_3 gnd vdd FILL
XFILL_87_DFFSR_218 gnd vdd FILL
XFILL_22_DFFSR_140 gnd vdd FILL
XFILL_87_DFFSR_229 gnd vdd FILL
XFILL_22_DFFSR_151 gnd vdd FILL
XFILL_22_DFFSR_162 gnd vdd FILL
XFILL_22_DFFSR_173 gnd vdd FILL
XFILL_3_INVX1_102 gnd vdd FILL
XFILL_22_DFFSR_184 gnd vdd FILL
XFILL_3_INVX1_113 gnd vdd FILL
XFILL_3_INVX1_124 gnd vdd FILL
XFILL_22_DFFSR_195 gnd vdd FILL
XFILL_1_NAND3X1_11 gnd vdd FILL
XFILL_3_INVX1_135 gnd vdd FILL
XFILL_3_INVX1_146 gnd vdd FILL
XFILL_1_NAND3X1_22 gnd vdd FILL
XFILL_3_INVX1_157 gnd vdd FILL
XFILL_1_NAND3X1_33 gnd vdd FILL
XFILL_3_INVX1_168 gnd vdd FILL
XFILL_26_DFFSR_150 gnd vdd FILL
XFILL_1_NAND3X1_44 gnd vdd FILL
XFILL_26_DFFSR_161 gnd vdd FILL
XFILL_1_NAND3X1_55 gnd vdd FILL
XFILL_1_NAND3X1_66 gnd vdd FILL
XFILL_26_DFFSR_172 gnd vdd FILL
XFILL_3_INVX1_179 gnd vdd FILL
XFILL_5_NAND2X1_13 gnd vdd FILL
XFILL_26_DFFSR_183 gnd vdd FILL
XFILL_5_NAND2X1_24 gnd vdd FILL
XFILL_7_INVX1_101 gnd vdd FILL
XFILL_1_NAND3X1_77 gnd vdd FILL
XFILL_7_INVX1_112 gnd vdd FILL
XFILL_5_NAND2X1_35 gnd vdd FILL
XFILL_7_INVX1_123 gnd vdd FILL
XFILL_1_NAND3X1_88 gnd vdd FILL
XFILL_26_DFFSR_194 gnd vdd FILL
XFILL_5_NAND2X1_46 gnd vdd FILL
XFILL_1_NAND3X1_99 gnd vdd FILL
XFILL_5_NAND2X1_57 gnd vdd FILL
XFILL_7_INVX1_134 gnd vdd FILL
XFILL_7_INVX1_145 gnd vdd FILL
XFILL_5_NAND2X1_68 gnd vdd FILL
XFILL_7_INVX1_156 gnd vdd FILL
XFILL_5_NAND2X1_79 gnd vdd FILL
XINVX1_170 INVX1_170/A gnd INVX1_170/Y vdd INVX1
XFILL_7_INVX1_167 gnd vdd FILL
XINVX1_181 INVX1_181/A gnd INVX1_181/Y vdd INVX1
XINVX1_192 DFFSR_94/Q gnd OAI21X1_6/A vdd INVX1
XFILL_7_INVX1_178 gnd vdd FILL
XFILL_7_INVX1_189 gnd vdd FILL
XFILL_22_NOR3X1_40 gnd vdd FILL
XFILL_22_NOR3X1_51 gnd vdd FILL
XFILL_1_OAI22X1_8 gnd vdd FILL
XFILL_72_DFFSR_240 gnd vdd FILL
XFILL_72_DFFSR_251 gnd vdd FILL
XFILL_72_DFFSR_262 gnd vdd FILL
XFILL_72_DFFSR_273 gnd vdd FILL
XFILL_26_NOR3X1_50 gnd vdd FILL
XFILL_11_NOR2X1_106 gnd vdd FILL
XFILL_5_OAI22X1_7 gnd vdd FILL
XFILL_11_NOR2X1_117 gnd vdd FILL
XFILL_11_NOR2X1_128 gnd vdd FILL
XFILL_76_DFFSR_250 gnd vdd FILL
XFILL_5_AOI22X1_11 gnd vdd FILL
XFILL_11_NOR2X1_139 gnd vdd FILL
XFILL_76_DFFSR_261 gnd vdd FILL
XFILL_52_3_0 gnd vdd FILL
XFILL_76_DFFSR_272 gnd vdd FILL
XFILL_31_CLKBUF1_2 gnd vdd FILL
XFILL_24_0_2 gnd vdd FILL
XFILL_50_DFFSR_208 gnd vdd FILL
XFILL_9_AOI21X1_13 gnd vdd FILL
XFILL_50_DFFSR_219 gnd vdd FILL
XFILL_9_OAI22X1_6 gnd vdd FILL
XFILL_9_AOI21X1_24 gnd vdd FILL
XFILL_9_AOI21X1_35 gnd vdd FILL
XFILL_9_AOI21X1_46 gnd vdd FILL
XFILL_35_CLKBUF1_1 gnd vdd FILL
XFILL_19_OAI22X1_15 gnd vdd FILL
XFILL_9_AOI21X1_57 gnd vdd FILL
XFILL_9_AOI21X1_68 gnd vdd FILL
XFILL_19_OAI22X1_26 gnd vdd FILL
XFILL_20_CLKBUF1_12 gnd vdd FILL
XFILL_9_AOI21X1_79 gnd vdd FILL
XFILL_20_CLKBUF1_23 gnd vdd FILL
XFILL_19_OAI22X1_37 gnd vdd FILL
XFILL_54_DFFSR_207 gnd vdd FILL
XFILL_20_CLKBUF1_34 gnd vdd FILL
XFILL_19_OAI22X1_48 gnd vdd FILL
XFILL_54_DFFSR_218 gnd vdd FILL
XFILL_54_DFFSR_229 gnd vdd FILL
XFILL_3_CLKBUF1_16 gnd vdd FILL
XFILL_3_CLKBUF1_27 gnd vdd FILL
XFILL_3_CLKBUF1_38 gnd vdd FILL
XFILL_81_DFFSR_107 gnd vdd FILL
XFILL_58_DFFSR_206 gnd vdd FILL
XFILL_81_DFFSR_118 gnd vdd FILL
XFILL_58_DFFSR_217 gnd vdd FILL
XFILL_58_DFFSR_228 gnd vdd FILL
XFILL_81_DFFSR_129 gnd vdd FILL
XFILL_58_DFFSR_239 gnd vdd FILL
XFILL_6_BUFX2_5 gnd vdd FILL
XFILL_85_DFFSR_106 gnd vdd FILL
XFILL_1_NOR2X1_101 gnd vdd FILL
XFILL_85_DFFSR_117 gnd vdd FILL
XFILL_1_NOR2X1_112 gnd vdd FILL
XFILL_12_OAI21X1_17 gnd vdd FILL
XFILL_1_NOR2X1_123 gnd vdd FILL
XFILL_85_DFFSR_128 gnd vdd FILL
XFILL_1_NOR2X1_134 gnd vdd FILL
XFILL_12_OAI21X1_28 gnd vdd FILL
XFILL_12_OAI21X1_39 gnd vdd FILL
XFILL_85_DFFSR_139 gnd vdd FILL
XFILL_1_NOR2X1_145 gnd vdd FILL
XFILL_7_1_2 gnd vdd FILL
XFILL_1_NOR2X1_156 gnd vdd FILL
XFILL_1_NOR2X1_167 gnd vdd FILL
XFILL_1_NOR2X1_178 gnd vdd FILL
XFILL_65_DFFSR_4 gnd vdd FILL
XFILL_8_BUFX4_13 gnd vdd FILL
XFILL_1_NOR2X1_189 gnd vdd FILL
XFILL_2_NAND3X1_9 gnd vdd FILL
XFILL_5_DFFSR_209 gnd vdd FILL
XFILL_8_BUFX4_24 gnd vdd FILL
XFILL_8_BUFX4_35 gnd vdd FILL
XFILL_4_OR2X2_1 gnd vdd FILL
XFILL_8_BUFX4_46 gnd vdd FILL
XFILL_11_NAND2X1_60 gnd vdd FILL
XFILL_8_BUFX4_57 gnd vdd FILL
XFILL_11_NAND2X1_71 gnd vdd FILL
XFILL_9_OAI22X1_10 gnd vdd FILL
XFILL_8_BUFX4_68 gnd vdd FILL
XFILL_11_NAND2X1_82 gnd vdd FILL
XFILL_9_OAI22X1_21 gnd vdd FILL
XFILL_9_OAI22X1_32 gnd vdd FILL
XFILL_8_BUFX4_79 gnd vdd FILL
XFILL_9_OAI22X1_43 gnd vdd FILL
XFILL_11_NAND2X1_93 gnd vdd FILL
XFILL_9_DFFSR_208 gnd vdd FILL
XFILL_6_NAND3X1_8 gnd vdd FILL
XFILL_9_DFFSR_219 gnd vdd FILL
XFILL_43_3_0 gnd vdd FILL
XFILL_15_0_2 gnd vdd FILL
XFILL_43_DFFSR_250 gnd vdd FILL
XNAND3X1_101 INVX1_83/A BUFX4_60/Y NOR2X1_44/Y gnd NAND3X1_102/A vdd NAND3X1
XFILL_43_DFFSR_261 gnd vdd FILL
XFILL_43_DFFSR_272 gnd vdd FILL
XFILL_1_MUX2X1_107 gnd vdd FILL
XNAND3X1_112 INVX1_172/A BUFX4_89/Y AND2X2_6/Y gnd NAND2X1_68/B vdd NAND3X1
XFILL_1_MUX2X1_118 gnd vdd FILL
XNAND3X1_123 DFFSR_21/Q BUFX4_8/Y NOR2X1_34/Y gnd NAND3X1_125/B vdd NAND3X1
XFILL_1_MUX2X1_129 gnd vdd FILL
XFILL_6_NOR2X1_201 gnd vdd FILL
XFILL_87_DFFSR_8 gnd vdd FILL
XFILL_70_DFFSR_150 gnd vdd FILL
XFILL_70_DFFSR_161 gnd vdd FILL
XFILL_15_AND2X2_1 gnd vdd FILL
XFILL_70_DFFSR_172 gnd vdd FILL
XFILL_47_DFFSR_260 gnd vdd FILL
XFILL_47_DFFSR_271 gnd vdd FILL
XFILL_2_OAI21X1_12 gnd vdd FILL
XFILL_70_DFFSR_183 gnd vdd FILL
XFILL_2_OAI21X1_23 gnd vdd FILL
XFILL_6_INVX2_5 gnd vdd FILL
XFILL_70_DFFSR_194 gnd vdd FILL
XFILL_21_DFFSR_207 gnd vdd FILL
XFILL_2_OAI21X1_34 gnd vdd FILL
XFILL_21_DFFSR_218 gnd vdd FILL
XFILL_2_OAI21X1_45 gnd vdd FILL
XFILL_21_DFFSR_229 gnd vdd FILL
XFILL_74_DFFSR_160 gnd vdd FILL
XFILL_74_DFFSR_171 gnd vdd FILL
XFILL_74_DFFSR_182 gnd vdd FILL
XFILL_74_DFFSR_193 gnd vdd FILL
XFILL_15_AOI21X1_60 gnd vdd FILL
XFILL_25_DFFSR_206 gnd vdd FILL
XFILL_15_AOI21X1_71 gnd vdd FILL
XFILL_25_DFFSR_217 gnd vdd FILL
XFILL_25_DFFSR_228 gnd vdd FILL
XFILL_4_INVX1_3 gnd vdd FILL
XFILL_12_BUFX4_40 gnd vdd FILL
XFILL_25_DFFSR_239 gnd vdd FILL
XFILL_21_DFFSR_19 gnd vdd FILL
XFILL_12_BUFX4_51 gnd vdd FILL
XFILL_78_DFFSR_170 gnd vdd FILL
XFILL_12_BUFX4_62 gnd vdd FILL
XFILL_12_BUFX4_73 gnd vdd FILL
XFILL_78_DFFSR_181 gnd vdd FILL
XFILL_12_BUFX4_84 gnd vdd FILL
XFILL_78_DFFSR_192 gnd vdd FILL
XFILL_52_DFFSR_106 gnd vdd FILL
XFILL_12_BUFX4_95 gnd vdd FILL
XFILL_29_DFFSR_205 gnd vdd FILL
XFILL_52_DFFSR_117 gnd vdd FILL
XFILL_29_DFFSR_216 gnd vdd FILL
XFILL_29_DFFSR_227 gnd vdd FILL
XFILL_52_DFFSR_128 gnd vdd FILL
XFILL_29_DFFSR_238 gnd vdd FILL
XFILL_61_DFFSR_18 gnd vdd FILL
XFILL_52_DFFSR_139 gnd vdd FILL
XFILL_29_DFFSR_249 gnd vdd FILL
XFILL_61_DFFSR_29 gnd vdd FILL
XFILL_56_DFFSR_105 gnd vdd FILL
XFILL_56_DFFSR_116 gnd vdd FILL
XFILL_56_DFFSR_127 gnd vdd FILL
XFILL_56_DFFSR_138 gnd vdd FILL
XFILL_56_DFFSR_149 gnd vdd FILL
XFILL_30_DFFSR_17 gnd vdd FILL
XFILL_34_3_0 gnd vdd FILL
XFILL_30_DFFSR_28 gnd vdd FILL
XFILL_30_DFFSR_39 gnd vdd FILL
XFILL_6_INVX1_30 gnd vdd FILL
XFILL_18_MUX2X1_110 gnd vdd FILL
XFILL_6_INVX1_41 gnd vdd FILL
XFILL_18_MUX2X1_121 gnd vdd FILL
XFILL_6_INVX1_52 gnd vdd FILL
XFILL_20_1 gnd vdd FILL
XFILL_18_MUX2X1_132 gnd vdd FILL
XFILL_6_INVX1_63 gnd vdd FILL
XFILL_6_INVX1_74 gnd vdd FILL
XFILL_18_MUX2X1_143 gnd vdd FILL
XFILL_10_DFFSR_250 gnd vdd FILL
XFILL_18_MUX2X1_154 gnd vdd FILL
XFILL_6_INVX1_85 gnd vdd FILL
XFILL_10_DFFSR_261 gnd vdd FILL
XFILL_18_MUX2X1_165 gnd vdd FILL
XFILL_3_DFFSR_108 gnd vdd FILL
XFILL_6_INVX1_96 gnd vdd FILL
XFILL_10_DFFSR_272 gnd vdd FILL
XFILL_70_DFFSR_16 gnd vdd FILL
XFILL_70_DFFSR_27 gnd vdd FILL
XFILL_3_DFFSR_119 gnd vdd FILL
XFILL_18_MUX2X1_176 gnd vdd FILL
XFILL_18_MUX2X1_187 gnd vdd FILL
XFILL_70_DFFSR_38 gnd vdd FILL
XFILL_70_DFFSR_49 gnd vdd FILL
XFILL_13_MUX2X1_6 gnd vdd FILL
XFILL_14_DFFSR_260 gnd vdd FILL
XDFFSR_110 INVX1_191/A DFFSR_78/CLK DFFSR_78/R vdd DFFSR_110/D gnd vdd DFFSR
XFILL_7_DFFSR_107 gnd vdd FILL
XFILL_14_DFFSR_271 gnd vdd FILL
XDFFSR_121 INVX1_175/A DFFSR_64/CLK DFFSR_2/R vdd DFFSR_121/D gnd vdd DFFSR
XDFFSR_132 INVX1_168/A DFFSR_55/CLK DFFSR_55/R vdd DFFSR_132/D gnd vdd DFFSR
XFILL_11_MUX2X1_16 gnd vdd FILL
XFILL_7_DFFSR_118 gnd vdd FILL
XDFFSR_143 INVX1_155/A DFFSR_72/CLK BUFX4_55/Y vdd DFFSR_143/D gnd vdd DFFSR
XFILL_7_DFFSR_129 gnd vdd FILL
XFILL_11_MUX2X1_27 gnd vdd FILL
XFILL_4_BUFX4_50 gnd vdd FILL
XDFFSR_154 INVX1_153/A DFFSR_81/CLK DFFSR_82/R vdd DFFSR_154/D gnd vdd DFFSR
XFILL_4_BUFX4_61 gnd vdd FILL
XFILL_11_MUX2X1_38 gnd vdd FILL
XFILL_2_AOI21X1_3 gnd vdd FILL
XDFFSR_165 INVX1_101/A CLKBUF1_6/Y DFFSR_56/R vdd MUX2X1_46/Y gnd vdd DFFSR
XFILL_11_MUX2X1_49 gnd vdd FILL
XBUFX4_6 BUFX4_8/A gnd BUFX4_6/Y vdd BUFX4
XFILL_4_BUFX4_72 gnd vdd FILL
XDFFSR_176 INVX1_24/A DFFSR_94/CLK DFFSR_98/R vdd DFFSR_176/D gnd vdd DFFSR
XFILL_4_BUFX4_83 gnd vdd FILL
XDFFSR_187 INVX1_133/A CLKBUF1_24/Y DFFSR_1/R vdd INVX1_131/A gnd vdd DFFSR
XFILL_41_DFFSR_160 gnd vdd FILL
XDFFSR_198 INVX1_98/A DFFSR_90/CLK BUFX4_32/Y vdd MUX2X1_85/Y gnd vdd DFFSR
XFILL_4_BUFX4_94 gnd vdd FILL
XFILL_41_DFFSR_171 gnd vdd FILL
XFILL_18_DFFSR_270 gnd vdd FILL
XFILL_15_MUX2X1_15 gnd vdd FILL
XFILL_41_DFFSR_182 gnd vdd FILL
XFILL_41_DFFSR_193 gnd vdd FILL
XFILL_15_MUX2X1_26 gnd vdd FILL
XFILL_15_MUX2X1_37 gnd vdd FILL
XFILL_6_AOI21X1_2 gnd vdd FILL
XFILL_15_MUX2X1_48 gnd vdd FILL
XFILL_15_MUX2X1_59 gnd vdd FILL
XFILL_45_DFFSR_170 gnd vdd FILL
XFILL_22_MUX2X1_4 gnd vdd FILL
XFILL_3_NOR3X1_19 gnd vdd FILL
XFILL_45_DFFSR_181 gnd vdd FILL
XFILL_19_MUX2X1_14 gnd vdd FILL
XFILL_19_MUX2X1_25 gnd vdd FILL
XFILL_45_DFFSR_192 gnd vdd FILL
XFILL_19_MUX2X1_36 gnd vdd FILL
XFILL_47_DFFSR_1 gnd vdd FILL
XFILL_19_MUX2X1_47 gnd vdd FILL
XNOR3X1_10 NOR3X1_10/A NOR3X1_46/B NOR3X1_46/C gnd NOR3X1_11/A vdd NOR3X1
XFILL_6_NOR2X1_7 gnd vdd FILL
XFILL_19_MUX2X1_58 gnd vdd FILL
XFILL_19_MUX2X1_69 gnd vdd FILL
XFILL_8_MUX2X1_160 gnd vdd FILL
XNOR3X1_21 INVX1_14/Y NOR3X1_5/B NOR3X1_5/C gnd NOR3X1_24/A vdd NOR3X1
XFILL_7_NOR3X1_18 gnd vdd FILL
XFILL_8_MUX2X1_171 gnd vdd FILL
XNOR3X1_32 NOR3X1_32/A NOR3X1_32/B NOR3X1_32/C gnd NOR3X1_32/Y vdd NOR3X1
XFILL_49_DFFSR_180 gnd vdd FILL
XFILL_8_MUX2X1_182 gnd vdd FILL
XNOR3X1_43 NOR3X1_43/A NOR3X1_43/B NOR3X1_43/C gnd NOR3X1_43/Y vdd NOR3X1
XFILL_7_NOR3X1_29 gnd vdd FILL
XFILL_49_DFFSR_191 gnd vdd FILL
XFILL_8_MUX2X1_193 gnd vdd FILL
XFILL_23_DFFSR_105 gnd vdd FILL
XFILL_23_DFFSR_116 gnd vdd FILL
XFILL_10_BUFX2_10 gnd vdd FILL
XFILL_23_DFFSR_127 gnd vdd FILL
XFILL_23_DFFSR_138 gnd vdd FILL
XFILL_23_DFFSR_149 gnd vdd FILL
XFILL_25_3_0 gnd vdd FILL
XFILL_0_3_0 gnd vdd FILL
XFILL_5_MUX2X1_5 gnd vdd FILL
XFILL_27_DFFSR_104 gnd vdd FILL
XFILL_27_DFFSR_115 gnd vdd FILL
XFILL_27_DFFSR_126 gnd vdd FILL
XFILL_27_DFFSR_137 gnd vdd FILL
XFILL_31_DFFSR_7 gnd vdd FILL
XFILL_27_DFFSR_148 gnd vdd FILL
XFILL_10_NAND3X1_13 gnd vdd FILL
XFILL_27_DFFSR_159 gnd vdd FILL
XFILL_10_NAND3X1_24 gnd vdd FILL
XFILL_10_NAND3X1_35 gnd vdd FILL
XFILL_10_NAND3X1_46 gnd vdd FILL
XFILL_69_DFFSR_5 gnd vdd FILL
XFILL_10_NAND3X1_57 gnd vdd FILL
XFILL_10_NAND3X1_68 gnd vdd FILL
XFILL_30_CLKBUF1_13 gnd vdd FILL
XFILL_30_CLKBUF1_24 gnd vdd FILL
XFILL_10_NAND3X1_79 gnd vdd FILL
XFILL_30_CLKBUF1_35 gnd vdd FILL
XFILL_39_DFFSR_50 gnd vdd FILL
XFILL_39_DFFSR_61 gnd vdd FILL
XFILL_39_DFFSR_72 gnd vdd FILL
XFILL_39_DFFSR_83 gnd vdd FILL
XFILL_23_NOR3X1_16 gnd vdd FILL
XFILL_39_DFFSR_94 gnd vdd FILL
XFILL_23_NOR3X1_27 gnd vdd FILL
XFILL_23_NOR3X1_38 gnd vdd FILL
XFILL_23_NOR3X1_49 gnd vdd FILL
XFILL_73_DFFSR_205 gnd vdd FILL
XFILL_0_DFFSR_13 gnd vdd FILL
XFILL_73_DFFSR_216 gnd vdd FILL
XFILL_0_DFFSR_24 gnd vdd FILL
XFILL_73_DFFSR_227 gnd vdd FILL
XFILL_73_DFFSR_238 gnd vdd FILL
XFILL_79_DFFSR_60 gnd vdd FILL
XFILL_10_NOR2X1_1 gnd vdd FILL
XFILL_0_DFFSR_35 gnd vdd FILL
XFILL_73_DFFSR_249 gnd vdd FILL
XFILL_79_DFFSR_71 gnd vdd FILL
XFILL_79_DFFSR_82 gnd vdd FILL
XFILL_0_DFFSR_46 gnd vdd FILL
XFILL_0_DFFSR_57 gnd vdd FILL
XFILL_79_DFFSR_93 gnd vdd FILL
XFILL_27_NOR3X1_15 gnd vdd FILL
XFILL_0_DFFSR_68 gnd vdd FILL
XFILL_27_NOR3X1_26 gnd vdd FILL
XFILL_0_DFFSR_79 gnd vdd FILL
XFILL_27_NOR3X1_37 gnd vdd FILL
XFILL_8_4_0 gnd vdd FILL
XFILL_27_NOR3X1_48 gnd vdd FILL
XFILL_77_DFFSR_204 gnd vdd FILL
XFILL_77_DFFSR_215 gnd vdd FILL
XFILL_77_DFFSR_226 gnd vdd FILL
XFILL_77_DFFSR_237 gnd vdd FILL
XFILL_77_DFFSR_248 gnd vdd FILL
XFILL_12_DFFSR_170 gnd vdd FILL
XFILL_19_NOR3X1_1 gnd vdd FILL
XFILL_1_CLKBUF1_2 gnd vdd FILL
XFILL_77_DFFSR_259 gnd vdd FILL
XFILL_12_DFFSR_181 gnd vdd FILL
XFILL_12_DFFSR_192 gnd vdd FILL
XFILL_48_DFFSR_70 gnd vdd FILL
XFILL_48_DFFSR_81 gnd vdd FILL
XFILL_48_DFFSR_92 gnd vdd FILL
XFILL_0_NAND3X1_30 gnd vdd FILL
XFILL_0_NAND3X1_41 gnd vdd FILL
XFILL_0_NAND3X1_52 gnd vdd FILL
XFILL_5_CLKBUF1_1 gnd vdd FILL
XFILL_4_NAND2X1_10 gnd vdd FILL
XFILL_0_NAND3X1_63 gnd vdd FILL
XFILL_16_DFFSR_180 gnd vdd FILL
XFILL_0_NAND3X1_74 gnd vdd FILL
XFILL_4_NAND2X1_21 gnd vdd FILL
XFILL_4_NAND2X1_32 gnd vdd FILL
XFILL_16_DFFSR_191 gnd vdd FILL
XFILL_0_NAND3X1_85 gnd vdd FILL
XFILL_4_NAND2X1_43 gnd vdd FILL
XFILL_0_NAND3X1_96 gnd vdd FILL
XFILL_16_3_0 gnd vdd FILL
XFILL_4_NAND2X1_54 gnd vdd FILL
XFILL_4_NAND2X1_65 gnd vdd FILL
XFILL_4_NAND2X1_76 gnd vdd FILL
XFILL_4_NAND2X1_87 gnd vdd FILL
XFILL_17_DFFSR_80 gnd vdd FILL
XFILL_17_DFFSR_91 gnd vdd FILL
XFILL_12_CLKBUF1_18 gnd vdd FILL
XFILL_12_CLKBUF1_29 gnd vdd FILL
XFILL_57_DFFSR_90 gnd vdd FILL
XFILL_62_DFFSR_270 gnd vdd FILL
XFILL_10_NOR2X1_103 gnd vdd FILL
XFILL_10_NOR2X1_114 gnd vdd FILL
XFILL_10_NOR2X1_125 gnd vdd FILL
XFILL_10_NOR2X1_136 gnd vdd FILL
XFILL_10_NOR2X1_147 gnd vdd FILL
XFILL_10_NOR2X1_158 gnd vdd FILL
XFILL_10_NOR2X1_169 gnd vdd FILL
XFILL_40_DFFSR_205 gnd vdd FILL
XFILL_8_AOI21X1_10 gnd vdd FILL
XFILL_40_DFFSR_216 gnd vdd FILL
XFILL_8_AOI21X1_21 gnd vdd FILL
XFILL_2_OAI21X1_6 gnd vdd FILL
XFILL_40_DFFSR_227 gnd vdd FILL
XFILL_8_AOI21X1_32 gnd vdd FILL
XFILL_40_DFFSR_238 gnd vdd FILL
XFILL_8_AOI21X1_43 gnd vdd FILL
XFILL_8_AOI21X1_54 gnd vdd FILL
XFILL_40_DFFSR_249 gnd vdd FILL
XFILL_18_OAI22X1_12 gnd vdd FILL
XFILL_18_OAI22X1_23 gnd vdd FILL
XNAND3X1_9 NOR2X1_96/Y NOR2X1_97/Y NOR3X1_38/Y gnd NOR3X1_43/C vdd NAND3X1
XFILL_8_AOI21X1_65 gnd vdd FILL
XFILL_18_OAI22X1_34 gnd vdd FILL
XFILL_8_AOI21X1_76 gnd vdd FILL
XFILL_44_DFFSR_204 gnd vdd FILL
XFILL_18_OAI22X1_45 gnd vdd FILL
XFILL_44_DFFSR_215 gnd vdd FILL
XFILL_3_NOR2X1_30 gnd vdd FILL
XFILL_6_OAI21X1_5 gnd vdd FILL
XFILL_3_NOR2X1_41 gnd vdd FILL
XFILL_44_DFFSR_226 gnd vdd FILL
XFILL_44_DFFSR_237 gnd vdd FILL
XFILL_66_2_0 gnd vdd FILL
XFILL_3_NOR2X1_52 gnd vdd FILL
XFILL_44_DFFSR_248 gnd vdd FILL
XFILL_3_NOR2X1_63 gnd vdd FILL
XFILL_13_BUFX4_18 gnd vdd FILL
XFILL_3_NOR2X1_74 gnd vdd FILL
XFILL_2_CLKBUF1_13 gnd vdd FILL
XFILL_44_DFFSR_259 gnd vdd FILL
XFILL_2_CLKBUF1_24 gnd vdd FILL
XFILL_13_BUFX4_29 gnd vdd FILL
XFILL_3_NOR2X1_85 gnd vdd FILL
XFILL_2_CLKBUF1_35 gnd vdd FILL
XFILL_71_DFFSR_104 gnd vdd FILL
XFILL_48_DFFSR_203 gnd vdd FILL
XFILL_3_NOR2X1_96 gnd vdd FILL
XFILL_10_MUX2X1_109 gnd vdd FILL
XFILL_71_DFFSR_115 gnd vdd FILL
XFILL_9_DFFSR_90 gnd vdd FILL
XFILL_71_DFFSR_126 gnd vdd FILL
XFILL_48_DFFSR_214 gnd vdd FILL
XFILL_48_DFFSR_225 gnd vdd FILL
XFILL_7_NOR2X1_40 gnd vdd FILL
XFILL_71_DFFSR_137 gnd vdd FILL
XFILL_7_NOR2X1_51 gnd vdd FILL
XFILL_48_DFFSR_236 gnd vdd FILL
XFILL_11_OAI22X1_2 gnd vdd FILL
XFILL_71_DFFSR_148 gnd vdd FILL
XFILL_48_DFFSR_247 gnd vdd FILL
XFILL_7_NOR2X1_62 gnd vdd FILL
XFILL_48_DFFSR_258 gnd vdd FILL
XFILL_71_DFFSR_159 gnd vdd FILL
XFILL_7_NOR2X1_73 gnd vdd FILL
XFILL_48_DFFSR_269 gnd vdd FILL
XFILL_7_NOR2X1_84 gnd vdd FILL
XFILL_7_NOR2X1_95 gnd vdd FILL
XFILL_75_DFFSR_103 gnd vdd FILL
XFILL_75_DFFSR_114 gnd vdd FILL
XFILL_11_OAI21X1_14 gnd vdd FILL
XFILL_50_6_1 gnd vdd FILL
XFILL_0_NOR2X1_120 gnd vdd FILL
XFILL_75_DFFSR_125 gnd vdd FILL
XFILL_75_DFFSR_136 gnd vdd FILL
XFILL_11_OAI21X1_25 gnd vdd FILL
XFILL_0_NOR2X1_131 gnd vdd FILL
XFILL_0_DFFSR_6 gnd vdd FILL
XFILL_11_OAI21X1_36 gnd vdd FILL
XFILL_15_OAI22X1_1 gnd vdd FILL
XFILL_11_OAI21X1_47 gnd vdd FILL
XFILL_75_DFFSR_147 gnd vdd FILL
XFILL_0_NOR2X1_142 gnd vdd FILL
XFILL_13_DFFSR_4 gnd vdd FILL
XFILL_75_DFFSR_158 gnd vdd FILL
XFILL_0_NOR2X1_153 gnd vdd FILL
XFILL_75_DFFSR_169 gnd vdd FILL
XFILL_0_NOR2X1_164 gnd vdd FILL
XFILL_70_DFFSR_5 gnd vdd FILL
XFILL_0_NOR2X1_175 gnd vdd FILL
XFILL_0_NOR2X1_186 gnd vdd FILL
XFILL_79_DFFSR_102 gnd vdd FILL
XFILL_0_NOR2X1_197 gnd vdd FILL
XFILL_79_DFFSR_113 gnd vdd FILL
XFILL_79_DFFSR_124 gnd vdd FILL
XFILL_79_DFFSR_135 gnd vdd FILL
XFILL_79_DFFSR_146 gnd vdd FILL
XFILL_79_DFFSR_157 gnd vdd FILL
XFILL_7_INVX1_19 gnd vdd FILL
XFILL_79_DFFSR_168 gnd vdd FILL
XFILL_10_NAND2X1_90 gnd vdd FILL
XFILL_79_DFFSR_179 gnd vdd FILL
XFILL_8_OAI22X1_40 gnd vdd FILL
XFILL_8_OAI22X1_51 gnd vdd FILL
XBUFX2_3 DFFSR_2/Q gnd dout[3] vdd BUFX2
XFILL_0_MUX2X1_104 gnd vdd FILL
XFILL_0_MUX2X1_115 gnd vdd FILL
XFILL_3_NAND2X1_7 gnd vdd FILL
XFILL_0_MUX2X1_126 gnd vdd FILL
XFILL_0_MUX2X1_137 gnd vdd FILL
XFILL_35_DFFSR_8 gnd vdd FILL
XFILL_0_MUX2X1_148 gnd vdd FILL
XFILL_5_BUFX4_17 gnd vdd FILL
XFILL_5_BUFX4_28 gnd vdd FILL
XFILL_0_MUX2X1_159 gnd vdd FILL
XFILL_5_BUFX4_39 gnd vdd FILL
XFILL_58_7_1 gnd vdd FILL
XFILL_60_DFFSR_180 gnd vdd FILL
XFILL_1_OAI21X1_20 gnd vdd FILL
XFILL_7_NAND2X1_6 gnd vdd FILL
XFILL_57_2_0 gnd vdd FILL
XFILL_1_OAI21X1_31 gnd vdd FILL
XFILL_60_DFFSR_191 gnd vdd FILL
XFILL_11_DFFSR_204 gnd vdd FILL
XFILL_11_DFFSR_215 gnd vdd FILL
XFILL_1_OAI21X1_42 gnd vdd FILL
XFILL_11_DFFSR_226 gnd vdd FILL
XFILL_11_DFFSR_237 gnd vdd FILL
XFILL_3_MUX2X1_70 gnd vdd FILL
XFILL_3_MUX2X1_81 gnd vdd FILL
XFILL_3_MUX2X1_92 gnd vdd FILL
XFILL_11_DFFSR_248 gnd vdd FILL
XFILL_11_DFFSR_259 gnd vdd FILL
XFILL_64_DFFSR_190 gnd vdd FILL
XFILL_12_NAND3X1_3 gnd vdd FILL
XFILL_15_DFFSR_203 gnd vdd FILL
XFILL_15_DFFSR_214 gnd vdd FILL
XFILL_15_DFFSR_225 gnd vdd FILL
XFILL_15_DFFSR_236 gnd vdd FILL
XFILL_7_MUX2X1_80 gnd vdd FILL
XFILL_15_DFFSR_247 gnd vdd FILL
XFILL_7_MUX2X1_91 gnd vdd FILL
XFILL_15_DFFSR_258 gnd vdd FILL
XFILL_15_DFFSR_269 gnd vdd FILL
XFILL_41_6_1 gnd vdd FILL
XFILL_19_DFFSR_202 gnd vdd FILL
XFILL_12_AND2X2_5 gnd vdd FILL
XFILL_42_DFFSR_103 gnd vdd FILL
XFILL_40_1_0 gnd vdd FILL
XFILL_42_DFFSR_114 gnd vdd FILL
XFILL_19_DFFSR_213 gnd vdd FILL
XFILL_42_DFFSR_125 gnd vdd FILL
XFILL_19_DFFSR_224 gnd vdd FILL
XFILL_42_DFFSR_136 gnd vdd FILL
XFILL_19_DFFSR_235 gnd vdd FILL
XINVX2_3 INVX2_3/A gnd INVX2_3/Y vdd INVX2
XFILL_19_DFFSR_246 gnd vdd FILL
XFILL_42_DFFSR_147 gnd vdd FILL
XFILL_42_DFFSR_158 gnd vdd FILL
XFILL_19_DFFSR_257 gnd vdd FILL
XFILL_42_DFFSR_169 gnd vdd FILL
XFILL_19_DFFSR_268 gnd vdd FILL
XFILL_46_DFFSR_102 gnd vdd FILL
XAOI21X1_3 BUFX4_99/Y AOI21X1_3/B AOI21X1_3/C gnd DFFSR_151/D vdd AOI21X1
XFILL_46_DFFSR_113 gnd vdd FILL
XFILL_46_DFFSR_124 gnd vdd FILL
XFILL_3_NAND3X1_18 gnd vdd FILL
XFILL_46_DFFSR_135 gnd vdd FILL
XFILL_3_NAND3X1_29 gnd vdd FILL
XFILL_46_DFFSR_146 gnd vdd FILL
XFILL_46_DFFSR_157 gnd vdd FILL
XFILL_46_DFFSR_168 gnd vdd FILL
XFILL_46_DFFSR_179 gnd vdd FILL
XMUX2X1_150 BUFX4_76/Y INVX1_194/Y NOR2X1_154/Y gnd DFFSR_96/D vdd MUX2X1
XMUX2X1_161 BUFX4_87/Y OAI21X1_5/A NOR2X1_162/Y gnd DFFSR_76/D vdd MUX2X1
XMUX2X1_172 BUFX4_76/Y INVX1_217/Y NOR2X1_165/Y gnd DFFSR_70/D vdd MUX2X1
XFILL_17_MUX2X1_140 gnd vdd FILL
XMUX2X1_183 BUFX4_80/Y OAI22X1_5/A NOR2X1_168/Y gnd DFFSR_54/D vdd MUX2X1
XFILL_12_AOI22X1_8 gnd vdd FILL
XMUX2X1_194 MUX2X1_6/B INVX1_15/Y MUX2X1_3/S gnd DFFSR_48/D vdd MUX2X1
XFILL_17_MUX2X1_151 gnd vdd FILL
XFILL_17_MUX2X1_162 gnd vdd FILL
XFILL_17_MUX2X1_173 gnd vdd FILL
XFILL_17_MUX2X1_184 gnd vdd FILL
XFILL_49_7_1 gnd vdd FILL
XFILL_48_2_0 gnd vdd FILL
XFILL_16_AOI22X1_7 gnd vdd FILL
XFILL_54_7 gnd vdd FILL
XINVX1_90 INVX1_90/A gnd INVX1_90/Y vdd INVX1
XBUFX2_10 BUFX2_10/A gnd dout[0] vdd BUFX2
XFILL_3_INVX1_12 gnd vdd FILL
XFILL_3_INVX1_23 gnd vdd FILL
XFILL_10_INVX8_2 gnd vdd FILL
XFILL_3_INVX1_34 gnd vdd FILL
XFILL_4_AND2X2_4 gnd vdd FILL
XFILL_3_INVX1_45 gnd vdd FILL
XFILL_3_INVX1_56 gnd vdd FILL
XFILL_3_INVX1_67 gnd vdd FILL
XFILL_3_INVX1_78 gnd vdd FILL
XFILL_31_DFFSR_190 gnd vdd FILL
XFILL_49_DFFSR_15 gnd vdd FILL
XFILL_3_INVX1_89 gnd vdd FILL
XFILL_49_DFFSR_26 gnd vdd FILL
XFILL_49_DFFSR_37 gnd vdd FILL
XFILL_49_DFFSR_48 gnd vdd FILL
XFILL_32_6_1 gnd vdd FILL
XFILL_49_DFFSR_59 gnd vdd FILL
XFILL_31_1_0 gnd vdd FILL
XFILL_1_BUFX4_10 gnd vdd FILL
XFILL_22_CLKBUF1_19 gnd vdd FILL
XFILL_1_BUFX4_21 gnd vdd FILL
XFILL_52_DFFSR_2 gnd vdd FILL
XFILL_1_BUFX4_32 gnd vdd FILL
XFILL_1_BUFX4_43 gnd vdd FILL
XFILL_1_BUFX4_54 gnd vdd FILL
XFILL_18_DFFSR_14 gnd vdd FILL
XFILL_1_BUFX4_65 gnd vdd FILL
XFILL_18_DFFSR_25 gnd vdd FILL
XFILL_18_DFFSR_36 gnd vdd FILL
XFILL_1_BUFX4_76 gnd vdd FILL
XFILL_18_DFFSR_47 gnd vdd FILL
XFILL_18_DFFSR_58 gnd vdd FILL
XFILL_7_MUX2X1_190 gnd vdd FILL
XFILL_1_BUFX4_87 gnd vdd FILL
XFILL_13_DFFSR_102 gnd vdd FILL
XFILL_1_BUFX4_98 gnd vdd FILL
XFILL_18_DFFSR_69 gnd vdd FILL
XFILL_13_DFFSR_113 gnd vdd FILL
XFILL_13_DFFSR_124 gnd vdd FILL
XFILL_58_DFFSR_13 gnd vdd FILL
XFILL_13_DFFSR_135 gnd vdd FILL
XFILL_13_DFFSR_146 gnd vdd FILL
XNOR2X1_1 INVX2_4/A INVX2_5/Y gnd NOR2X1_1/Y vdd NOR2X1
XFILL_13_DFFSR_157 gnd vdd FILL
XFILL_58_DFFSR_24 gnd vdd FILL
XFILL_58_DFFSR_35 gnd vdd FILL
XFILL_13_DFFSR_168 gnd vdd FILL
XFILL_13_DFFSR_179 gnd vdd FILL
XFILL_58_DFFSR_46 gnd vdd FILL
XFILL_58_DFFSR_57 gnd vdd FILL
XFILL_17_DFFSR_101 gnd vdd FILL
XFILL_58_DFFSR_68 gnd vdd FILL
XFILL_17_DFFSR_112 gnd vdd FILL
XFILL_58_DFFSR_79 gnd vdd FILL
XFILL_3_NOR2X1_108 gnd vdd FILL
XFILL_17_DFFSR_123 gnd vdd FILL
XFILL_17_DFFSR_134 gnd vdd FILL
XFILL_3_NOR2X1_119 gnd vdd FILL
XFILL_4_DFFSR_7 gnd vdd FILL
XFILL_17_DFFSR_145 gnd vdd FILL
XFILL_17_DFFSR_5 gnd vdd FILL
XFILL_17_DFFSR_156 gnd vdd FILL
XFILL_17_DFFSR_167 gnd vdd FILL
XFILL_17_DFFSR_178 gnd vdd FILL
XFILL_74_DFFSR_6 gnd vdd FILL
XFILL_27_DFFSR_12 gnd vdd FILL
XFILL_17_DFFSR_189 gnd vdd FILL
XFILL_27_DFFSR_23 gnd vdd FILL
XFILL_39_2_0 gnd vdd FILL
XFILL_27_DFFSR_34 gnd vdd FILL
XFILL_27_DFFSR_45 gnd vdd FILL
XFILL_27_DFFSR_56 gnd vdd FILL
XFILL_27_DFFSR_67 gnd vdd FILL
XFILL_27_DFFSR_78 gnd vdd FILL
XFILL_2_BUFX4_105 gnd vdd FILL
XFILL_27_DFFSR_89 gnd vdd FILL
XFILL_13_NOR3X1_13 gnd vdd FILL
XFILL_67_DFFSR_11 gnd vdd FILL
XFILL_13_NOR3X1_24 gnd vdd FILL
XFILL_67_DFFSR_22 gnd vdd FILL
XFILL_13_NOR3X1_35 gnd vdd FILL
XFILL_67_DFFSR_33 gnd vdd FILL
XFILL_63_DFFSR_202 gnd vdd FILL
XFILL_13_NOR3X1_46 gnd vdd FILL
XFILL_67_DFFSR_44 gnd vdd FILL
XFILL_2_MUX2X1_9 gnd vdd FILL
XFILL_67_DFFSR_55 gnd vdd FILL
XFILL_63_DFFSR_213 gnd vdd FILL
XFILL_67_DFFSR_66 gnd vdd FILL
XFILL_63_DFFSR_224 gnd vdd FILL
XFILL_67_DFFSR_77 gnd vdd FILL
XFILL_63_DFFSR_235 gnd vdd FILL
XFILL_6_BUFX4_104 gnd vdd FILL
XFILL_67_DFFSR_88 gnd vdd FILL
XFILL_63_DFFSR_246 gnd vdd FILL
XFILL_17_NOR3X1_12 gnd vdd FILL
XFILL_67_DFFSR_99 gnd vdd FILL
XFILL_23_6_1 gnd vdd FILL
XFILL_63_DFFSR_257 gnd vdd FILL
XFILL_63_DFFSR_268 gnd vdd FILL
XFILL_17_NOR3X1_23 gnd vdd FILL
XFILL_17_NOR3X1_34 gnd vdd FILL
XFILL_67_DFFSR_201 gnd vdd FILL
XFILL_22_1_0 gnd vdd FILL
XFILL_17_NOR3X1_45 gnd vdd FILL
XFILL_39_DFFSR_9 gnd vdd FILL
XFILL_67_DFFSR_212 gnd vdd FILL
XFILL_36_DFFSR_10 gnd vdd FILL
XFILL_36_DFFSR_21 gnd vdd FILL
XFILL_67_DFFSR_223 gnd vdd FILL
XFILL_67_DFFSR_234 gnd vdd FILL
XFILL_0_OAI22X1_17 gnd vdd FILL
XFILL_36_DFFSR_32 gnd vdd FILL
XFILL_36_DFFSR_43 gnd vdd FILL
XFILL_67_DFFSR_245 gnd vdd FILL
XFILL_0_OAI22X1_28 gnd vdd FILL
XFILL_67_DFFSR_256 gnd vdd FILL
XFILL_0_OAI22X1_39 gnd vdd FILL
XFILL_36_DFFSR_54 gnd vdd FILL
XFILL_67_DFFSR_267 gnd vdd FILL
XFILL_22_CLKBUF1_8 gnd vdd FILL
XFILL_36_DFFSR_65 gnd vdd FILL
XFILL_36_DFFSR_76 gnd vdd FILL
XFILL_13_AOI22X1_10 gnd vdd FILL
XFILL_4_OAI21X1_19 gnd vdd FILL
XAOI21X1_11 BUFX4_98/Y AOI21X1_9/B NOR2X1_147/Y gnd DFFSR_106/D vdd AOI21X1
XFILL_36_DFFSR_87 gnd vdd FILL
XFILL_0_NOR2X1_18 gnd vdd FILL
XFILL_36_DFFSR_98 gnd vdd FILL
XAOI21X1_22 MUX2X1_66/A MUX2X1_14/S NOR2X1_176/Y gnd DFFSR_36/D vdd AOI21X1
XFILL_0_NOR2X1_29 gnd vdd FILL
XAOI21X1_33 BUFX4_99/Y NOR2X1_190/B NOR2X1_190/Y gnd DFFSR_22/D vdd AOI21X1
XAOI21X1_44 BUFX4_97/Y MUX2X1_22/S NOR2X1_205/Y gnd DFFSR_5/D vdd AOI21X1
XFILL_76_DFFSR_20 gnd vdd FILL
XFILL_76_DFFSR_31 gnd vdd FILL
XFILL_76_DFFSR_42 gnd vdd FILL
XAOI21X1_55 BUFX4_97/Y NOR2X1_16/B NOR2X1_16/Y gnd DFFSR_261/D vdd AOI21X1
XAOI21X1_66 DFFSR_148/Q NOR2X1_43/Y NOR2X1_47/Y gnd NAND3X1_50/B vdd AOI21X1
XFILL_76_DFFSR_53 gnd vdd FILL
XAOI21X1_77 NOR2X1_21/A NAND2X1_92/Y INVX1_141/Y gnd NOR3X1_48/B vdd AOI21X1
XFILL_26_CLKBUF1_7 gnd vdd FILL
XFILL_76_DFFSR_64 gnd vdd FILL
XFILL_76_DFFSR_75 gnd vdd FILL
XFILL_3_NAND2X1_40 gnd vdd FILL
XFILL_76_DFFSR_86 gnd vdd FILL
XFILL_3_NAND2X1_51 gnd vdd FILL
XOAI21X1_6 OAI21X1_6/A OAI21X1_6/B OAI21X1_6/C gnd OAI21X1_6/Y vdd OAI21X1
XFILL_3_NAND2X1_62 gnd vdd FILL
XFILL_76_DFFSR_97 gnd vdd FILL
XFILL_4_NOR2X1_17 gnd vdd FILL
XFILL_4_NOR2X1_28 gnd vdd FILL
XFILL_3_NAND2X1_73 gnd vdd FILL
XFILL_4_NOR2X1_39 gnd vdd FILL
XFILL_11_BUFX4_5 gnd vdd FILL
XFILL_3_NAND2X1_84 gnd vdd FILL
XFILL_3_NAND2X1_95 gnd vdd FILL
XFILL_45_DFFSR_30 gnd vdd FILL
XFILL_45_DFFSR_41 gnd vdd FILL
XFILL_11_CLKBUF1_15 gnd vdd FILL
XFILL_16_NOR3X1_5 gnd vdd FILL
XFILL_11_CLKBUF1_26 gnd vdd FILL
XFILL_45_DFFSR_52 gnd vdd FILL
XFILL_8_NOR2X1_16 gnd vdd FILL
XFILL_45_DFFSR_63 gnd vdd FILL
XFILL_8_NOR2X1_27 gnd vdd FILL
XFILL_11_CLKBUF1_37 gnd vdd FILL
XFILL_8_NOR2X1_38 gnd vdd FILL
XFILL_6_7_1 gnd vdd FILL
XFILL_45_DFFSR_74 gnd vdd FILL
XFILL_8_NOR2X1_49 gnd vdd FILL
XFILL_45_DFFSR_85 gnd vdd FILL
XFILL_45_DFFSR_96 gnd vdd FILL
XFILL_5_2_0 gnd vdd FILL
XFILL_85_DFFSR_40 gnd vdd FILL
XFILL_85_DFFSR_51 gnd vdd FILL
XFILL_85_DFFSR_62 gnd vdd FILL
XFILL_85_DFFSR_73 gnd vdd FILL
XFILL_85_DFFSR_84 gnd vdd FILL
XFILL_14_DFFSR_40 gnd vdd FILL
XFILL_85_DFFSR_95 gnd vdd FILL
XFILL_14_DFFSR_51 gnd vdd FILL
XFILL_14_DFFSR_62 gnd vdd FILL
XFILL_14_DFFSR_73 gnd vdd FILL
XFILL_14_DFFSR_84 gnd vdd FILL
XFILL_14_DFFSR_95 gnd vdd FILL
XFILL_30_DFFSR_202 gnd vdd FILL
XFILL_30_DFFSR_213 gnd vdd FILL
XFILL_25_NOR3X1_3 gnd vdd FILL
XFILL_14_6_1 gnd vdd FILL
XFILL_30_DFFSR_224 gnd vdd FILL
XFILL_30_DFFSR_235 gnd vdd FILL
XOAI22X1_30 INVX1_1/Y OAI22X1_4/B INVX1_24/Y OAI22X1_4/D gnd NOR2X1_93/B vdd OAI22X1
XOAI22X1_41 MUX2X1_95/A OAI22X1_7/D MUX2X1_99/A NOR2X1_60/B gnd OAI22X1_41/Y vdd OAI22X1
XFILL_7_AOI21X1_40 gnd vdd FILL
XFILL_13_1_0 gnd vdd FILL
XFILL_30_DFFSR_246 gnd vdd FILL
XFILL_54_DFFSR_50 gnd vdd FILL
XFILL_7_AOI21X1_51 gnd vdd FILL
XFILL_54_DFFSR_61 gnd vdd FILL
XFILL_7_AOI21X1_62 gnd vdd FILL
XFILL_30_DFFSR_257 gnd vdd FILL
XFILL_54_DFFSR_72 gnd vdd FILL
XFILL_54_DFFSR_83 gnd vdd FILL
XFILL_30_DFFSR_268 gnd vdd FILL
XFILL_17_OAI22X1_20 gnd vdd FILL
XFILL_17_OAI22X1_31 gnd vdd FILL
XFILL_7_AOI21X1_73 gnd vdd FILL
XFILL_34_DFFSR_201 gnd vdd FILL
XFILL_17_OAI22X1_42 gnd vdd FILL
XFILL_54_DFFSR_94 gnd vdd FILL
XFILL_34_DFFSR_212 gnd vdd FILL
XFILL_34_DFFSR_223 gnd vdd FILL
XFILL_34_DFFSR_234 gnd vdd FILL
XFILL_34_DFFSR_245 gnd vdd FILL
XFILL_1_CLKBUF1_10 gnd vdd FILL
XFILL_34_DFFSR_256 gnd vdd FILL
XFILL_1_CLKBUF1_21 gnd vdd FILL
XFILL_34_DFFSR_267 gnd vdd FILL
XFILL_0_MUX2X1_14 gnd vdd FILL
XFILL_1_CLKBUF1_32 gnd vdd FILL
XFILL_0_MUX2X1_25 gnd vdd FILL
XFILL_61_DFFSR_101 gnd vdd FILL
XFILL_38_DFFSR_200 gnd vdd FILL
XFILL_0_MUX2X1_36 gnd vdd FILL
XFILL_38_DFFSR_211 gnd vdd FILL
XFILL_23_DFFSR_60 gnd vdd FILL
XFILL_61_DFFSR_112 gnd vdd FILL
XFILL_0_MUX2X1_47 gnd vdd FILL
XFILL_23_DFFSR_71 gnd vdd FILL
XFILL_61_DFFSR_123 gnd vdd FILL
XFILL_23_DFFSR_82 gnd vdd FILL
XFILL_61_DFFSR_134 gnd vdd FILL
XFILL_38_DFFSR_222 gnd vdd FILL
XFILL_0_MUX2X1_58 gnd vdd FILL
XFILL_14_INVX8_3 gnd vdd FILL
XFILL_0_MUX2X1_69 gnd vdd FILL
XFILL_23_DFFSR_93 gnd vdd FILL
XFILL_38_DFFSR_233 gnd vdd FILL
XFILL_61_DFFSR_145 gnd vdd FILL
XFILL_38_DFFSR_244 gnd vdd FILL
XFILL_8_NOR3X1_4 gnd vdd FILL
XFILL_61_DFFSR_156 gnd vdd FILL
XFILL_38_DFFSR_255 gnd vdd FILL
XFILL_61_DFFSR_167 gnd vdd FILL
XFILL_38_DFFSR_266 gnd vdd FILL
XFILL_61_DFFSR_178 gnd vdd FILL
XFILL_4_MUX2X1_13 gnd vdd FILL
XFILL_4_MUX2X1_24 gnd vdd FILL
XFILL_65_DFFSR_100 gnd vdd FILL
XFILL_4_MUX2X1_35 gnd vdd FILL
XFILL_61_DFFSR_189 gnd vdd FILL
XFILL_10_OAI21X1_11 gnd vdd FILL
XFILL_65_DFFSR_111 gnd vdd FILL
XFILL_4_MUX2X1_46 gnd vdd FILL
XFILL_63_DFFSR_70 gnd vdd FILL
XFILL_65_DFFSR_122 gnd vdd FILL
XFILL_65_DFFSR_133 gnd vdd FILL
XFILL_63_DFFSR_81 gnd vdd FILL
XFILL_4_MUX2X1_57 gnd vdd FILL
XFILL_10_OAI21X1_22 gnd vdd FILL
XFILL_63_DFFSR_92 gnd vdd FILL
XFILL_65_DFFSR_144 gnd vdd FILL
XFILL_4_MUX2X1_68 gnd vdd FILL
XFILL_10_OAI21X1_33 gnd vdd FILL
XFILL_4_MUX2X1_79 gnd vdd FILL
XFILL_10_OAI21X1_44 gnd vdd FILL
XFILL_65_DFFSR_155 gnd vdd FILL
XFILL_3_3 gnd vdd FILL
XFILL_65_DFFSR_166 gnd vdd FILL
XFILL_65_DFFSR_177 gnd vdd FILL
XFILL_8_MUX2X1_12 gnd vdd FILL
XFILL_8_MUX2X1_23 gnd vdd FILL
XFILL_65_DFFSR_188 gnd vdd FILL
XFILL_8_MUX2X1_34 gnd vdd FILL
XFILL_56_DFFSR_3 gnd vdd FILL
XFILL_8_MUX2X1_45 gnd vdd FILL
XFILL_69_DFFSR_110 gnd vdd FILL
XFILL_65_DFFSR_199 gnd vdd FILL
XFILL_69_DFFSR_121 gnd vdd FILL
XFILL_6_DFFSR_50 gnd vdd FILL
XFILL_69_DFFSR_132 gnd vdd FILL
XFILL_8_MUX2X1_56 gnd vdd FILL
XFILL_6_DFFSR_61 gnd vdd FILL
XFILL_69_DFFSR_143 gnd vdd FILL
XFILL_6_DFFSR_72 gnd vdd FILL
XFILL_8_MUX2X1_67 gnd vdd FILL
XFILL_6_DFFSR_83 gnd vdd FILL
XFILL_8_MUX2X1_78 gnd vdd FILL
XFILL_69_DFFSR_154 gnd vdd FILL
XFILL_6_DFFSR_94 gnd vdd FILL
XFILL_8_MUX2X1_89 gnd vdd FILL
XFILL_69_DFFSR_165 gnd vdd FILL
XFILL_32_DFFSR_80 gnd vdd FILL
XFILL_69_DFFSR_176 gnd vdd FILL
XFILL_64_5_1 gnd vdd FILL
XFILL_32_DFFSR_91 gnd vdd FILL
XFILL_69_DFFSR_187 gnd vdd FILL
XFILL_69_DFFSR_198 gnd vdd FILL
XFILL_45_3 gnd vdd FILL
XFILL_63_0_0 gnd vdd FILL
XFILL_38_2 gnd vdd FILL
XFILL_72_DFFSR_90 gnd vdd FILL
XFILL_20_MUX2X1_11 gnd vdd FILL
XFILL_20_MUX2X1_22 gnd vdd FILL
XFILL_40_DFFSR_9 gnd vdd FILL
XFILL_20_MUX2X1_33 gnd vdd FILL
XFILL_8_DFFSR_8 gnd vdd FILL
XFILL_20_MUX2X1_44 gnd vdd FILL
XFILL_20_MUX2X1_55 gnd vdd FILL
XFILL_20_MUX2X1_66 gnd vdd FILL
XFILL_20_MUX2X1_77 gnd vdd FILL
XFILL_20_MUX2X1_88 gnd vdd FILL
XFILL_78_DFFSR_7 gnd vdd FILL
XFILL_20_MUX2X1_99 gnd vdd FILL
XFILL_0_OAI21X1_50 gnd vdd FILL
XFILL_32_DFFSR_100 gnd vdd FILL
XFILL_32_DFFSR_111 gnd vdd FILL
XFILL_32_DFFSR_122 gnd vdd FILL
XFILL_32_DFFSR_133 gnd vdd FILL
XFILL_32_DFFSR_144 gnd vdd FILL
XFILL_32_DFFSR_155 gnd vdd FILL
XFILL_32_DFFSR_166 gnd vdd FILL
XFILL_32_DFFSR_177 gnd vdd FILL
XFILL_1_DFFSR_190 gnd vdd FILL
XFILL_32_DFFSR_188 gnd vdd FILL
XFILL_36_DFFSR_110 gnd vdd FILL
XFILL_32_DFFSR_199 gnd vdd FILL
XFILL_2_NAND3X1_15 gnd vdd FILL
XFILL_36_DFFSR_121 gnd vdd FILL
XFILL_36_DFFSR_132 gnd vdd FILL
XFILL_2_NAND3X1_26 gnd vdd FILL
XFILL_55_5_1 gnd vdd FILL
XFILL_36_DFFSR_143 gnd vdd FILL
XFILL_2_NAND3X1_37 gnd vdd FILL
XFILL_36_DFFSR_154 gnd vdd FILL
XFILL_2_NAND3X1_48 gnd vdd FILL
XFILL_54_0_0 gnd vdd FILL
XFILL_2_NAND3X1_59 gnd vdd FILL
XFILL_36_DFFSR_165 gnd vdd FILL
XFILL_36_DFFSR_176 gnd vdd FILL
XFILL_6_NAND2X1_17 gnd vdd FILL
XFILL_6_NAND2X1_28 gnd vdd FILL
XFILL_36_DFFSR_187 gnd vdd FILL
XFILL_36_DFFSR_198 gnd vdd FILL
XFILL_6_NAND2X1_39 gnd vdd FILL
XFILL_2_BUFX4_8 gnd vdd FILL
XFILL_15_BUFX4_6 gnd vdd FILL
XFILL_16_MUX2X1_170 gnd vdd FILL
XFILL_16_MUX2X1_181 gnd vdd FILL
XFILL_82_DFFSR_200 gnd vdd FILL
XFILL_16_MUX2X1_192 gnd vdd FILL
XFILL_82_DFFSR_211 gnd vdd FILL
XFILL_82_DFFSR_222 gnd vdd FILL
XFILL_82_DFFSR_233 gnd vdd FILL
XFILL_82_DFFSR_244 gnd vdd FILL
XFILL_82_DFFSR_255 gnd vdd FILL
XFILL_82_DFFSR_266 gnd vdd FILL
XFILL_86_DFFSR_210 gnd vdd FILL
XFILL_86_DFFSR_221 gnd vdd FILL
XFILL_13_AOI21X1_6 gnd vdd FILL
XFILL_86_DFFSR_232 gnd vdd FILL
XFILL_86_DFFSR_243 gnd vdd FILL
XFILL_86_DFFSR_254 gnd vdd FILL
XFILL_86_DFFSR_265 gnd vdd FILL
XFILL_11_BUFX2_2 gnd vdd FILL
XFILL_2_INVX1_160 gnd vdd FILL
XFILL_2_INVX1_171 gnd vdd FILL
XFILL_2_INVX1_182 gnd vdd FILL
XFILL_2_INVX1_193 gnd vdd FILL
XFILL_21_CLKBUF1_16 gnd vdd FILL
XFILL_21_CLKBUF1_27 gnd vdd FILL
XFILL_21_CLKBUF1_38 gnd vdd FILL
XBUFX4_105 BUFX4_8/A gnd NAND3X1_7/B vdd BUFX4
XFILL_6_INVX1_170 gnd vdd FILL
XFILL_0_INVX1_16 gnd vdd FILL
XFILL_6_INVX1_181 gnd vdd FILL
XFILL_0_INVX1_27 gnd vdd FILL
XFILL_6_INVX1_192 gnd vdd FILL
XFILL_0_INVX1_38 gnd vdd FILL
XFILL_46_5_1 gnd vdd FILL
XFILL_1_AND2X2_8 gnd vdd FILL
XFILL_0_INVX1_49 gnd vdd FILL
XFILL_45_0_0 gnd vdd FILL
XFILL_18_INVX8_4 gnd vdd FILL
XFILL_46_DFFSR_19 gnd vdd FILL
XFILL_31_9 gnd vdd FILL
XFILL_24_8 gnd vdd FILL
XFILL_2_NOR2X1_105 gnd vdd FILL
XFILL_2_NOR2X1_116 gnd vdd FILL
XFILL_2_NOR2X1_127 gnd vdd FILL
XFILL_86_DFFSR_18 gnd vdd FILL
XFILL_86_DFFSR_29 gnd vdd FILL
XFILL_2_NOR2X1_138 gnd vdd FILL
XFILL_22_DFFSR_6 gnd vdd FILL
XFILL_2_NOR2X1_149 gnd vdd FILL
XFILL_15_DFFSR_18 gnd vdd FILL
XFILL_15_DFFSR_29 gnd vdd FILL
XFILL_55_DFFSR_17 gnd vdd FILL
XFILL_55_DFFSR_28 gnd vdd FILL
XFILL_55_DFFSR_39 gnd vdd FILL
XFILL_53_DFFSR_210 gnd vdd FILL
XFILL_53_DFFSR_221 gnd vdd FILL
XFILL_53_DFFSR_232 gnd vdd FILL
XFILL_53_DFFSR_243 gnd vdd FILL
XFILL_53_DFFSR_254 gnd vdd FILL
XFILL_53_DFFSR_265 gnd vdd FILL
XFILL_9_NAND3X1_90 gnd vdd FILL
XFILL_24_DFFSR_16 gnd vdd FILL
XFILL_80_DFFSR_110 gnd vdd FILL
XFILL_7_NOR2X1_205 gnd vdd FILL
XFILL_24_DFFSR_27 gnd vdd FILL
XFILL_80_DFFSR_121 gnd vdd FILL
XFILL_80_DFFSR_132 gnd vdd FILL
XFILL_57_DFFSR_220 gnd vdd FILL
XFILL_15_BUFX4_70 gnd vdd FILL
XFILL_24_DFFSR_38 gnd vdd FILL
XFILL_57_DFFSR_231 gnd vdd FILL
XFILL_80_DFFSR_143 gnd vdd FILL
XFILL_57_DFFSR_242 gnd vdd FILL
XFILL_24_DFFSR_49 gnd vdd FILL
XFILL_80_DFFSR_154 gnd vdd FILL
XFILL_15_BUFX4_81 gnd vdd FILL
XFILL_57_DFFSR_253 gnd vdd FILL
XFILL_15_BUFX4_92 gnd vdd FILL
XFILL_80_DFFSR_165 gnd vdd FILL
XFILL_57_DFFSR_264 gnd vdd FILL
XFILL_80_DFFSR_176 gnd vdd FILL
XFILL_12_CLKBUF1_5 gnd vdd FILL
XFILL_0_DFFSR_202 gnd vdd FILL
XFILL_57_DFFSR_275 gnd vdd FILL
XFILL_3_OAI21X1_16 gnd vdd FILL
XFILL_80_DFFSR_187 gnd vdd FILL
XFILL_3_OAI21X1_27 gnd vdd FILL
XFILL_0_DFFSR_213 gnd vdd FILL
XFILL_80_DFFSR_198 gnd vdd FILL
XFILL_3_OAI21X1_38 gnd vdd FILL
XFILL_64_DFFSR_15 gnd vdd FILL
XFILL_50_1 gnd vdd FILL
XFILL_84_DFFSR_120 gnd vdd FILL
XFILL_64_DFFSR_26 gnd vdd FILL
XFILL_0_DFFSR_224 gnd vdd FILL
XFILL_84_DFFSR_131 gnd vdd FILL
XFILL_0_DFFSR_235 gnd vdd FILL
XFILL_3_OAI21X1_49 gnd vdd FILL
XFILL_64_DFFSR_37 gnd vdd FILL
XFILL_84_DFFSR_142 gnd vdd FILL
XFILL_37_5_1 gnd vdd FILL
XFILL_0_DFFSR_246 gnd vdd FILL
XFILL_64_DFFSR_48 gnd vdd FILL
XFILL_84_DFFSR_153 gnd vdd FILL
XFILL_0_DFFSR_257 gnd vdd FILL
XFILL_64_DFFSR_59 gnd vdd FILL
XFILL_0_DFFSR_268 gnd vdd FILL
XFILL_36_0_0 gnd vdd FILL
XFILL_84_DFFSR_164 gnd vdd FILL
XFILL_84_DFFSR_175 gnd vdd FILL
XFILL_16_CLKBUF1_4 gnd vdd FILL
XFILL_4_DFFSR_201 gnd vdd FILL
XFILL_84_DFFSR_186 gnd vdd FILL
XFILL_84_DFFSR_197 gnd vdd FILL
XFILL_4_DFFSR_212 gnd vdd FILL
XFILL_1_NAND3X1_1 gnd vdd FILL
XFILL_4_DFFSR_223 gnd vdd FILL
XFILL_4_DFFSR_234 gnd vdd FILL
XFILL_7_DFFSR_17 gnd vdd FILL
XFILL_2_NAND2X1_70 gnd vdd FILL
XFILL_2_NAND2X1_81 gnd vdd FILL
XFILL_7_DFFSR_28 gnd vdd FILL
XFILL_4_DFFSR_245 gnd vdd FILL
XFILL_2_NAND2X1_92 gnd vdd FILL
XFILL_4_DFFSR_256 gnd vdd FILL
XFILL_33_DFFSR_14 gnd vdd FILL
XFILL_7_DFFSR_39 gnd vdd FILL
XFILL_4_DFFSR_267 gnd vdd FILL
XFILL_33_DFFSR_25 gnd vdd FILL
XFILL_33_DFFSR_36 gnd vdd FILL
XFILL_8_DFFSR_200 gnd vdd FILL
XFILL_33_DFFSR_47 gnd vdd FILL
XFILL_10_CLKBUF1_12 gnd vdd FILL
XFILL_8_DFFSR_211 gnd vdd FILL
XFILL_10_CLKBUF1_23 gnd vdd FILL
XFILL_33_DFFSR_58 gnd vdd FILL
XFILL_39_DFFSR_209 gnd vdd FILL
XFILL_10_CLKBUF1_34 gnd vdd FILL
XFILL_8_DFFSR_222 gnd vdd FILL
XFILL_33_DFFSR_69 gnd vdd FILL
XFILL_8_DFFSR_233 gnd vdd FILL
XFILL_8_DFFSR_244 gnd vdd FILL
XFILL_20_4_1 gnd vdd FILL
XFILL_8_DFFSR_255 gnd vdd FILL
XFILL_73_DFFSR_13 gnd vdd FILL
XFILL_8_DFFSR_266 gnd vdd FILL
XFILL_73_DFFSR_24 gnd vdd FILL
XFILL_73_DFFSR_35 gnd vdd FILL
XFILL_73_DFFSR_46 gnd vdd FILL
XFILL_73_DFFSR_57 gnd vdd FILL
XFILL_16_MUX2X1_3 gnd vdd FILL
XFILL_66_DFFSR_109 gnd vdd FILL
XFILL_73_DFFSR_68 gnd vdd FILL
XFILL_73_DFFSR_79 gnd vdd FILL
XFILL_6_BUFX4_9 gnd vdd FILL
XFILL_42_DFFSR_12 gnd vdd FILL
XFILL_7_BUFX4_80 gnd vdd FILL
XFILL_42_DFFSR_23 gnd vdd FILL
XFILL_19_MUX2X1_103 gnd vdd FILL
XFILL_20_DFFSR_210 gnd vdd FILL
XFILL_42_DFFSR_34 gnd vdd FILL
XFILL_10_NOR2X1_12 gnd vdd FILL
XFILL_19_MUX2X1_114 gnd vdd FILL
XFILL_7_BUFX4_91 gnd vdd FILL
XFILL_13_NOR3X1_9 gnd vdd FILL
XFILL_20_DFFSR_221 gnd vdd FILL
XFILL_42_DFFSR_45 gnd vdd FILL
XFILL_10_NOR2X1_23 gnd vdd FILL
XFILL_1_AOI22X1_6 gnd vdd FILL
XFILL_42_DFFSR_56 gnd vdd FILL
XFILL_19_MUX2X1_125 gnd vdd FILL
XFILL_20_DFFSR_232 gnd vdd FILL
XFILL_10_NOR2X1_34 gnd vdd FILL
XFILL_20_DFFSR_243 gnd vdd FILL
XFILL_13_OAI21X1_9 gnd vdd FILL
XFILL_42_DFFSR_67 gnd vdd FILL
XFILL_19_MUX2X1_136 gnd vdd FILL
XFILL_10_NOR2X1_45 gnd vdd FILL
XFILL_20_DFFSR_254 gnd vdd FILL
XFILL_19_MUX2X1_147 gnd vdd FILL
XFILL_10_NOR2X1_56 gnd vdd FILL
XFILL_42_DFFSR_78 gnd vdd FILL
XFILL_42_DFFSR_89 gnd vdd FILL
XFILL_6_AOI21X1_70 gnd vdd FILL
XFILL_19_MUX2X1_158 gnd vdd FILL
XFILL_10_NOR2X1_67 gnd vdd FILL
XFILL_20_DFFSR_265 gnd vdd FILL
XFILL_10_NOR2X1_78 gnd vdd FILL
XFILL_1_INVX1_205 gnd vdd FILL
XFILL_82_DFFSR_11 gnd vdd FILL
XFILL_19_MUX2X1_169 gnd vdd FILL
XFILL_6_AOI21X1_81 gnd vdd FILL
XFILL_82_DFFSR_22 gnd vdd FILL
XFILL_10_NOR2X1_89 gnd vdd FILL
XFILL_16_OAI22X1_50 gnd vdd FILL
XFILL_1_INVX1_216 gnd vdd FILL
XFILL_1_INVX1_227 gnd vdd FILL
XFILL_82_DFFSR_33 gnd vdd FILL
XFILL_5_AOI22X1_5 gnd vdd FILL
XFILL_24_DFFSR_220 gnd vdd FILL
XFILL_82_DFFSR_44 gnd vdd FILL
XFILL_82_DFFSR_55 gnd vdd FILL
XFILL_11_DFFSR_11 gnd vdd FILL
XFILL_24_DFFSR_231 gnd vdd FILL
XFILL_24_DFFSR_242 gnd vdd FILL
XFILL_11_DFFSR_22 gnd vdd FILL
XFILL_82_DFFSR_66 gnd vdd FILL
XFILL_82_DFFSR_77 gnd vdd FILL
XFILL_24_DFFSR_253 gnd vdd FILL
XFILL_24_DFFSR_264 gnd vdd FILL
XFILL_11_DFFSR_33 gnd vdd FILL
XFILL_82_DFFSR_88 gnd vdd FILL
XFILL_11_DFFSR_44 gnd vdd FILL
XFILL_24_DFFSR_275 gnd vdd FILL
XFILL_11_DFFSR_55 gnd vdd FILL
XFILL_82_DFFSR_99 gnd vdd FILL
XFILL_5_INVX1_204 gnd vdd FILL
XFILL_28_5_1 gnd vdd FILL
XFILL_11_DFFSR_66 gnd vdd FILL
XFILL_3_5_1 gnd vdd FILL
XFILL_9_NOR2X1_180 gnd vdd FILL
XFILL_0_CLKBUF1_40 gnd vdd FILL
XFILL_11_DFFSR_77 gnd vdd FILL
XFILL_5_INVX1_215 gnd vdd FILL
XFILL_9_NOR2X1_191 gnd vdd FILL
XFILL_9_NOR2X1_4 gnd vdd FILL
XFILL_51_DFFSR_120 gnd vdd FILL
XFILL_5_INVX1_226 gnd vdd FILL
XFILL_27_0_0 gnd vdd FILL
XFILL_51_DFFSR_131 gnd vdd FILL
XFILL_2_0_0 gnd vdd FILL
XFILL_11_DFFSR_88 gnd vdd FILL
XFILL_9_AOI22X1_4 gnd vdd FILL
XFILL_51_DFFSR_142 gnd vdd FILL
XFILL_11_DFFSR_99 gnd vdd FILL
XFILL_28_DFFSR_230 gnd vdd FILL
XFILL_51_DFFSR_10 gnd vdd FILL
XFILL_51_DFFSR_21 gnd vdd FILL
XFILL_28_DFFSR_241 gnd vdd FILL
XFILL_51_DFFSR_153 gnd vdd FILL
XFILL_28_DFFSR_252 gnd vdd FILL
XFILL_51_DFFSR_32 gnd vdd FILL
XFILL_2_BUFX2_5 gnd vdd FILL
XFILL_22_NOR3X1_7 gnd vdd FILL
XFILL_28_DFFSR_263 gnd vdd FILL
XFILL_51_DFFSR_164 gnd vdd FILL
XFILL_51_DFFSR_43 gnd vdd FILL
XFILL_51_DFFSR_175 gnd vdd FILL
XFILL_28_DFFSR_274 gnd vdd FILL
XFILL_51_DFFSR_186 gnd vdd FILL
XFILL_51_DFFSR_54 gnd vdd FILL
XFILL_51_DFFSR_65 gnd vdd FILL
XFILL_51_DFFSR_76 gnd vdd FILL
XFILL_51_DFFSR_197 gnd vdd FILL
XFILL_51_DFFSR_87 gnd vdd FILL
XFILL_55_DFFSR_130 gnd vdd FILL
XFILL_51_DFFSR_98 gnd vdd FILL
XFILL_55_DFFSR_141 gnd vdd FILL
XFILL_8_MUX2X1_2 gnd vdd FILL
XFILL_55_DFFSR_152 gnd vdd FILL
XFILL_55_DFFSR_163 gnd vdd FILL
XFILL_55_DFFSR_174 gnd vdd FILL
XFILL_11_4_1 gnd vdd FILL
XFILL_55_DFFSR_185 gnd vdd FILL
XFILL_61_DFFSR_4 gnd vdd FILL
XFILL_20_DFFSR_20 gnd vdd FILL
XFILL_55_DFFSR_196 gnd vdd FILL
XFILL_9_MUX2X1_120 gnd vdd FILL
XFILL_20_DFFSR_31 gnd vdd FILL
XFILL_20_DFFSR_42 gnd vdd FILL
XFILL_9_MUX2X1_131 gnd vdd FILL
XFILL_59_DFFSR_140 gnd vdd FILL
XFILL_0_OR2X2_1 gnd vdd FILL
XFILL_9_MUX2X1_142 gnd vdd FILL
XFILL_20_DFFSR_53 gnd vdd FILL
XFILL_9_MUX2X1_153 gnd vdd FILL
XFILL_59_DFFSR_151 gnd vdd FILL
XFILL_20_DFFSR_64 gnd vdd FILL
XFILL_9_MUX2X1_164 gnd vdd FILL
XFILL_20_DFFSR_75 gnd vdd FILL
XFILL_59_DFFSR_162 gnd vdd FILL
XFILL_20_DFFSR_86 gnd vdd FILL
XFILL_9_MUX2X1_175 gnd vdd FILL
XFILL_59_DFFSR_173 gnd vdd FILL
XFILL_20_DFFSR_97 gnd vdd FILL
XFILL_59_DFFSR_184 gnd vdd FILL
XFILL_5_NOR3X1_8 gnd vdd FILL
XFILL_9_MUX2X1_186 gnd vdd FILL
XFILL_2_DFFSR_100 gnd vdd FILL
XFILL_59_DFFSR_195 gnd vdd FILL
XFILL_2_DFFSR_111 gnd vdd FILL
XFILL_33_DFFSR_109 gnd vdd FILL
XFILL_60_DFFSR_30 gnd vdd FILL
XFILL_2_DFFSR_122 gnd vdd FILL
XFILL_2_DFFSR_133 gnd vdd FILL
XFILL_60_DFFSR_41 gnd vdd FILL
XFILL_31_NOR3X1_5 gnd vdd FILL
XFILL_2_DFFSR_144 gnd vdd FILL
XFILL_60_DFFSR_52 gnd vdd FILL
XFILL_60_DFFSR_63 gnd vdd FILL
XFILL_2_DFFSR_155 gnd vdd FILL
XFILL_60_DFFSR_74 gnd vdd FILL
XFILL_2_DFFSR_166 gnd vdd FILL
XFILL_2_DFFSR_177 gnd vdd FILL
XFILL_60_DFFSR_85 gnd vdd FILL
XFILL_60_DFFSR_96 gnd vdd FILL
XFILL_2_DFFSR_188 gnd vdd FILL
XFILL_6_DFFSR_110 gnd vdd FILL
XFILL_2_DFFSR_199 gnd vdd FILL
XFILL_37_DFFSR_108 gnd vdd FILL
XFILL_6_DFFSR_121 gnd vdd FILL
XFILL_3_DFFSR_10 gnd vdd FILL
XFILL_3_DFFSR_21 gnd vdd FILL
XFILL_6_DFFSR_132 gnd vdd FILL
XFILL_10_MUX2X1_30 gnd vdd FILL
XFILL_37_DFFSR_119 gnd vdd FILL
XFILL_6_DFFSR_143 gnd vdd FILL
XFILL_10_MUX2X1_41 gnd vdd FILL
XFILL_3_DFFSR_32 gnd vdd FILL
XFILL_3_DFFSR_43 gnd vdd FILL
XFILL_6_DFFSR_154 gnd vdd FILL
XFILL_10_MUX2X1_52 gnd vdd FILL
XFILL_26_DFFSR_7 gnd vdd FILL
XFILL_11_NAND3X1_17 gnd vdd FILL
XFILL_6_DFFSR_165 gnd vdd FILL
XFILL_10_MUX2X1_63 gnd vdd FILL
XFILL_3_DFFSR_54 gnd vdd FILL
XFILL_83_DFFSR_8 gnd vdd FILL
XFILL_3_DFFSR_65 gnd vdd FILL
XFILL_11_NAND3X1_28 gnd vdd FILL
XFILL_10_MUX2X1_74 gnd vdd FILL
XFILL_6_DFFSR_176 gnd vdd FILL
XFILL_3_DFFSR_76 gnd vdd FILL
XFILL_10_MUX2X1_85 gnd vdd FILL
XFILL_6_DFFSR_187 gnd vdd FILL
XFILL_11_NAND3X1_39 gnd vdd FILL
XFILL_10_MUX2X1_96 gnd vdd FILL
XFILL_6_DFFSR_198 gnd vdd FILL
XFILL_3_DFFSR_87 gnd vdd FILL
XFILL_3_DFFSR_98 gnd vdd FILL
XFILL_2_INVX2_5 gnd vdd FILL
XFILL_31_CLKBUF1_17 gnd vdd FILL
XFILL_31_CLKBUF1_28 gnd vdd FILL
XFILL_14_MUX2X1_40 gnd vdd FILL
XFILL_14_MUX2X1_51 gnd vdd FILL
XFILL_31_CLKBUF1_39 gnd vdd FILL
XFILL_19_5_1 gnd vdd FILL
XFILL_14_MUX2X1_62 gnd vdd FILL
XFILL_14_MUX2X1_73 gnd vdd FILL
XFILL_2_NOR3X1_11 gnd vdd FILL
XFILL_14_MUX2X1_84 gnd vdd FILL
XFILL_18_0_0 gnd vdd FILL
XFILL_2_NOR3X1_22 gnd vdd FILL
XFILL_14_MUX2X1_95 gnd vdd FILL
XFILL_2_NOR3X1_33 gnd vdd FILL
XFILL_2_NOR3X1_44 gnd vdd FILL
XFILL_83_DFFSR_209 gnd vdd FILL
XFILL_18_MUX2X1_50 gnd vdd FILL
XFILL_18_MUX2X1_61 gnd vdd FILL
XFILL_0_INVX1_3 gnd vdd FILL
XFILL_61_3_1 gnd vdd FILL
XFILL_6_NOR3X1_10 gnd vdd FILL
XFILL_18_MUX2X1_72 gnd vdd FILL
XFILL_18_MUX2X1_83 gnd vdd FILL
XFILL_6_NOR3X1_21 gnd vdd FILL
XFILL_18_MUX2X1_94 gnd vdd FILL
XFILL_6_NOR3X1_32 gnd vdd FILL
XFILL_22_5 gnd vdd FILL
XFILL_6_NOR3X1_43 gnd vdd FILL
XFILL_87_DFFSR_208 gnd vdd FILL
XFILL_22_DFFSR_130 gnd vdd FILL
XFILL_87_DFFSR_219 gnd vdd FILL
XFILL_15_4 gnd vdd FILL
XFILL_22_DFFSR_141 gnd vdd FILL
XFILL_22_DFFSR_152 gnd vdd FILL
XFILL_22_DFFSR_163 gnd vdd FILL
XFILL_22_DFFSR_174 gnd vdd FILL
XFILL_3_INVX1_103 gnd vdd FILL
XFILL_22_DFFSR_185 gnd vdd FILL
XFILL_3_INVX1_114 gnd vdd FILL
XFILL_22_DFFSR_196 gnd vdd FILL
XFILL_3_INVX1_125 gnd vdd FILL
XFILL_1_NAND3X1_12 gnd vdd FILL
XFILL_3_INVX1_136 gnd vdd FILL
XFILL_1_NAND3X1_23 gnd vdd FILL
XFILL_3_INVX1_147 gnd vdd FILL
XFILL_26_DFFSR_140 gnd vdd FILL
XFILL_1_NAND3X1_34 gnd vdd FILL
XFILL_26_DFFSR_151 gnd vdd FILL
XFILL_3_INVX1_158 gnd vdd FILL
XFILL_3_INVX1_169 gnd vdd FILL
XFILL_1_NAND3X1_45 gnd vdd FILL
XFILL_26_DFFSR_162 gnd vdd FILL
XFILL_5_NAND2X1_14 gnd vdd FILL
XFILL_1_NAND3X1_56 gnd vdd FILL
XFILL_7_INVX1_102 gnd vdd FILL
XFILL_26_DFFSR_173 gnd vdd FILL
XFILL_1_NAND3X1_67 gnd vdd FILL
XFILL_26_DFFSR_184 gnd vdd FILL
XFILL_1_NAND3X1_78 gnd vdd FILL
XFILL_5_NAND2X1_25 gnd vdd FILL
XFILL_1_NAND3X1_89 gnd vdd FILL
XFILL_5_NAND2X1_36 gnd vdd FILL
XFILL_7_INVX1_113 gnd vdd FILL
XFILL_26_DFFSR_195 gnd vdd FILL
XFILL_7_INVX1_124 gnd vdd FILL
XFILL_5_NAND2X1_47 gnd vdd FILL
XFILL_5_NAND2X1_58 gnd vdd FILL
XFILL_7_INVX1_135 gnd vdd FILL
XFILL_7_INVX1_146 gnd vdd FILL
XINVX1_160 NOR2X1_7/A gnd INVX1_160/Y vdd INVX1
XFILL_5_NAND2X1_69 gnd vdd FILL
XFILL_7_INVX1_157 gnd vdd FILL
XINVX1_171 INVX1_171/A gnd INVX1_171/Y vdd INVX1
XFILL_7_INVX1_168 gnd vdd FILL
XINVX1_182 INVX1_182/A gnd INVX1_182/Y vdd INVX1
XINVX1_193 DFFSR_95/Q gnd INVX1_193/Y vdd INVX1
XFILL_7_INVX1_179 gnd vdd FILL
XFILL_22_NOR3X1_30 gnd vdd FILL
XFILL_22_NOR3X1_41 gnd vdd FILL
XFILL_22_NOR3X1_52 gnd vdd FILL
XFILL_72_DFFSR_230 gnd vdd FILL
XFILL_1_OAI22X1_9 gnd vdd FILL
XFILL_72_DFFSR_241 gnd vdd FILL
XFILL_72_DFFSR_252 gnd vdd FILL
XFILL_72_DFFSR_263 gnd vdd FILL
XFILL_72_DFFSR_274 gnd vdd FILL
XFILL_26_NOR3X1_40 gnd vdd FILL
XFILL_26_NOR3X1_51 gnd vdd FILL
XFILL_5_OAI22X1_8 gnd vdd FILL
XFILL_11_NOR2X1_107 gnd vdd FILL
XFILL_11_NOR2X1_118 gnd vdd FILL
XFILL_11_NOR2X1_129 gnd vdd FILL
XFILL_1_NOR3X1_1 gnd vdd FILL
XFILL_76_DFFSR_240 gnd vdd FILL
XFILL_76_DFFSR_251 gnd vdd FILL
XFILL_76_DFFSR_262 gnd vdd FILL
XFILL_31_CLKBUF1_3 gnd vdd FILL
XFILL_76_DFFSR_273 gnd vdd FILL
XFILL_52_3_1 gnd vdd FILL
XFILL_9_AOI21X1_14 gnd vdd FILL
XFILL_50_DFFSR_209 gnd vdd FILL
XFILL_9_OAI22X1_7 gnd vdd FILL
XFILL_9_AOI21X1_25 gnd vdd FILL
XFILL_9_AOI21X1_36 gnd vdd FILL
XFILL_9_AOI21X1_47 gnd vdd FILL
XFILL_9_AOI21X1_58 gnd vdd FILL
XFILL_9_AOI21X1_69 gnd vdd FILL
XFILL_19_OAI22X1_16 gnd vdd FILL
XFILL_35_CLKBUF1_2 gnd vdd FILL
XFILL_19_OAI22X1_27 gnd vdd FILL
XFILL_20_CLKBUF1_13 gnd vdd FILL
XFILL_19_OAI22X1_38 gnd vdd FILL
XFILL_54_DFFSR_208 gnd vdd FILL
XFILL_20_CLKBUF1_24 gnd vdd FILL
XFILL_19_OAI22X1_49 gnd vdd FILL
XFILL_20_CLKBUF1_35 gnd vdd FILL
XFILL_54_DFFSR_219 gnd vdd FILL
XFILL_43_DFFSR_1 gnd vdd FILL
XFILL_3_CLKBUF1_17 gnd vdd FILL
XFILL_3_CLKBUF1_28 gnd vdd FILL
XFILL_3_CLKBUF1_39 gnd vdd FILL
XFILL_58_DFFSR_207 gnd vdd FILL
XFILL_81_DFFSR_108 gnd vdd FILL
XFILL_81_DFFSR_119 gnd vdd FILL
XFILL_58_DFFSR_218 gnd vdd FILL
XFILL_58_DFFSR_229 gnd vdd FILL
XFILL_6_BUFX2_6 gnd vdd FILL
XFILL_1_NOR2X1_102 gnd vdd FILL
XFILL_85_DFFSR_107 gnd vdd FILL
XFILL_1_NOR2X1_113 gnd vdd FILL
XFILL_12_OAI21X1_18 gnd vdd FILL
XFILL_85_DFFSR_118 gnd vdd FILL
XFILL_1_NOR2X1_124 gnd vdd FILL
XFILL_85_DFFSR_129 gnd vdd FILL
XFILL_12_OAI21X1_29 gnd vdd FILL
XFILL_1_NOR2X1_135 gnd vdd FILL
XFILL_1_NOR2X1_146 gnd vdd FILL
XFILL_1_NOR2X1_157 gnd vdd FILL
XFILL_1_NOR2X1_168 gnd vdd FILL
XFILL_65_DFFSR_5 gnd vdd FILL
XFILL_1_NOR2X1_179 gnd vdd FILL
XFILL_8_BUFX4_14 gnd vdd FILL
XFILL_8_BUFX4_25 gnd vdd FILL
XFILL_11_NAND2X1_50 gnd vdd FILL
XFILL_8_BUFX4_36 gnd vdd FILL
XFILL_8_BUFX4_47 gnd vdd FILL
XFILL_9_OAI22X1_11 gnd vdd FILL
XFILL_11_NAND2X1_61 gnd vdd FILL
XFILL_8_BUFX4_58 gnd vdd FILL
XFILL_8_BUFX4_69 gnd vdd FILL
XFILL_11_NAND2X1_72 gnd vdd FILL
XFILL_9_OAI22X1_22 gnd vdd FILL
XFILL_11_NAND2X1_83 gnd vdd FILL
XFILL_11_NAND2X1_94 gnd vdd FILL
XFILL_9_OAI22X1_33 gnd vdd FILL
XFILL_9_OAI22X1_44 gnd vdd FILL
XFILL_9_DFFSR_209 gnd vdd FILL
XFILL_6_NAND3X1_9 gnd vdd FILL
XFILL_43_3_1 gnd vdd FILL
XFILL_43_DFFSR_240 gnd vdd FILL
XFILL_43_DFFSR_251 gnd vdd FILL
XNAND3X1_102 NAND3X1_102/A NAND3X1_98/Y NAND3X1_99/Y gnd NOR3X1_28/B vdd NAND3X1
XFILL_43_DFFSR_262 gnd vdd FILL
XFILL_1_MUX2X1_108 gnd vdd FILL
XNAND3X1_113 INVX1_153/A BUFX4_91/Y NOR2X1_44/Y gnd NAND2X1_69/A vdd NAND3X1
XFILL_43_DFFSR_273 gnd vdd FILL
XFILL_1_MUX2X1_119 gnd vdd FILL
XNAND3X1_124 DFFSR_17/Q BUFX4_8/Y NOR2X1_36/Y gnd NAND3X1_125/C vdd NAND3X1
XFILL_6_NOR2X1_202 gnd vdd FILL
XFILL_70_DFFSR_140 gnd vdd FILL
XFILL_87_DFFSR_9 gnd vdd FILL
XFILL_70_DFFSR_151 gnd vdd FILL
XFILL_47_DFFSR_250 gnd vdd FILL
XFILL_70_DFFSR_162 gnd vdd FILL
XFILL_15_AND2X2_2 gnd vdd FILL
XFILL_47_DFFSR_261 gnd vdd FILL
XFILL_47_DFFSR_272 gnd vdd FILL
XFILL_70_DFFSR_173 gnd vdd FILL
XFILL_70_DFFSR_184 gnd vdd FILL
XFILL_2_OAI21X1_13 gnd vdd FILL
XFILL_2_OAI21X1_24 gnd vdd FILL
XFILL_70_DFFSR_195 gnd vdd FILL
XFILL_21_DFFSR_208 gnd vdd FILL
XFILL_2_OAI21X1_35 gnd vdd FILL
XFILL_2_OAI21X1_46 gnd vdd FILL
XFILL_21_DFFSR_219 gnd vdd FILL
XFILL_74_DFFSR_150 gnd vdd FILL
XFILL_74_DFFSR_161 gnd vdd FILL
XFILL_74_DFFSR_172 gnd vdd FILL
XFILL_15_AOI21X1_50 gnd vdd FILL
XFILL_74_DFFSR_183 gnd vdd FILL
XFILL_74_DFFSR_194 gnd vdd FILL
XFILL_25_DFFSR_207 gnd vdd FILL
XFILL_15_AOI21X1_61 gnd vdd FILL
XFILL_15_AOI21X1_72 gnd vdd FILL
XFILL_4_INVX1_4 gnd vdd FILL
XFILL_25_DFFSR_218 gnd vdd FILL
XFILL_12_BUFX4_30 gnd vdd FILL
XFILL_25_DFFSR_229 gnd vdd FILL
XFILL_12_BUFX4_41 gnd vdd FILL
XFILL_78_DFFSR_160 gnd vdd FILL
XFILL_12_BUFX4_52 gnd vdd FILL
XFILL_12_BUFX4_63 gnd vdd FILL
XFILL_78_DFFSR_171 gnd vdd FILL
XFILL_12_BUFX4_74 gnd vdd FILL
XFILL_78_DFFSR_182 gnd vdd FILL
XFILL_12_BUFX4_85 gnd vdd FILL
XFILL_78_DFFSR_193 gnd vdd FILL
XFILL_29_DFFSR_206 gnd vdd FILL
XFILL_52_DFFSR_107 gnd vdd FILL
XFILL_12_BUFX4_96 gnd vdd FILL
XFILL_29_DFFSR_217 gnd vdd FILL
XFILL_52_DFFSR_118 gnd vdd FILL
XFILL_52_DFFSR_129 gnd vdd FILL
XFILL_6_10 gnd vdd FILL
XFILL_29_DFFSR_228 gnd vdd FILL
XFILL_61_DFFSR_19 gnd vdd FILL
XFILL_29_DFFSR_239 gnd vdd FILL
XFILL_56_DFFSR_106 gnd vdd FILL
XFILL_56_DFFSR_117 gnd vdd FILL
XFILL_56_DFFSR_128 gnd vdd FILL
XFILL_56_DFFSR_139 gnd vdd FILL
XFILL_30_DFFSR_18 gnd vdd FILL
XFILL_34_3_1 gnd vdd FILL
XFILL_30_DFFSR_29 gnd vdd FILL
XFILL_6_INVX1_20 gnd vdd FILL
XFILL_18_MUX2X1_100 gnd vdd FILL
XFILL_6_INVX1_31 gnd vdd FILL
XFILL_6_INVX1_42 gnd vdd FILL
XFILL_18_MUX2X1_111 gnd vdd FILL
XFILL_7_AND2X2_1 gnd vdd FILL
XFILL_18_MUX2X1_122 gnd vdd FILL
XFILL_6_INVX1_53 gnd vdd FILL
XFILL_6_INVX1_64 gnd vdd FILL
XFILL_10_DFFSR_240 gnd vdd FILL
XFILL_20_2 gnd vdd FILL
XFILL_18_MUX2X1_133 gnd vdd FILL
XFILL_18_MUX2X1_144 gnd vdd FILL
XFILL_10_DFFSR_251 gnd vdd FILL
XFILL_6_INVX1_75 gnd vdd FILL
XFILL_6_INVX1_86 gnd vdd FILL
XFILL_18_MUX2X1_155 gnd vdd FILL
XFILL_10_DFFSR_262 gnd vdd FILL
XFILL_6_INVX1_97 gnd vdd FILL
XFILL_3_DFFSR_109 gnd vdd FILL
XFILL_70_DFFSR_17 gnd vdd FILL
XFILL_10_DFFSR_273 gnd vdd FILL
XFILL_13_1 gnd vdd FILL
XFILL_18_MUX2X1_166 gnd vdd FILL
XFILL_70_DFFSR_28 gnd vdd FILL
XFILL_18_MUX2X1_177 gnd vdd FILL
XFILL_18_MUX2X1_188 gnd vdd FILL
XFILL_70_DFFSR_39 gnd vdd FILL
XFILL_13_MUX2X1_7 gnd vdd FILL
XDFFSR_100 DFFSR_100/Q DFFSR_93/CLK DFFSR_93/R vdd DFFSR_100/D gnd vdd DFFSR
XFILL_14_DFFSR_250 gnd vdd FILL
XDFFSR_111 INVX1_183/A CLKBUF1_31/Y DFFSR_64/R vdd DFFSR_111/D gnd vdd DFFSR
XFILL_14_DFFSR_261 gnd vdd FILL
XFILL_14_DFFSR_272 gnd vdd FILL
XFILL_7_DFFSR_108 gnd vdd FILL
XDFFSR_122 INVX1_176/A CLKBUF1_34/Y BUFX4_23/Y vdd DFFSR_122/D gnd vdd DFFSR
XDFFSR_133 INVX1_169/A DFFSR_58/CLK DFFSR_91/R vdd DFFSR_133/D gnd vdd DFFSR
XFILL_7_DFFSR_119 gnd vdd FILL
XFILL_11_MUX2X1_17 gnd vdd FILL
XDFFSR_144 INVX1_156/A DFFSR_72/CLK BUFX4_55/Y vdd DFFSR_144/D gnd vdd DFFSR
XFILL_4_BUFX4_40 gnd vdd FILL
XFILL_11_MUX2X1_28 gnd vdd FILL
XFILL_4_BUFX4_51 gnd vdd FILL
XDFFSR_155 INVX1_154/A CLKBUF1_31/Y DFFSR_53/R vdd DFFSR_155/D gnd vdd DFFSR
XFILL_11_MUX2X1_39 gnd vdd FILL
XDFFSR_166 INVX1_135/A DFFSR_52/CLK DFFSR_42/R vdd MUX2X1_57/Y gnd vdd DFFSR
XFILL_4_BUFX4_62 gnd vdd FILL
XFILL_2_AOI21X1_4 gnd vdd FILL
XFILL_4_BUFX4_73 gnd vdd FILL
XBUFX4_7 BUFX4_8/A gnd BUFX4_7/Y vdd BUFX4
XFILL_4_BUFX4_84 gnd vdd FILL
XDFFSR_177 INVX1_35/A DFFSR_70/CLK BUFX4_55/Y vdd MUX2X1_2/Y gnd vdd DFFSR
XFILL_41_DFFSR_150 gnd vdd FILL
XDFFSR_188 INVX1_132/A DFFSR_6/CLK DFFSR_6/R vdd INVX1_130/A gnd vdd DFFSR
XFILL_41_DFFSR_161 gnd vdd FILL
XFILL_4_BUFX4_95 gnd vdd FILL
XFILL_18_DFFSR_260 gnd vdd FILL
XDFFSR_199 INVX2_3/A DFFSR_1/CLK DFFSR_1/R vdd DFFSR_199/D gnd vdd DFFSR
XFILL_18_DFFSR_271 gnd vdd FILL
XFILL_41_DFFSR_172 gnd vdd FILL
XFILL_41_DFFSR_183 gnd vdd FILL
XFILL_15_MUX2X1_16 gnd vdd FILL
XFILL_41_DFFSR_194 gnd vdd FILL
XFILL_15_MUX2X1_27 gnd vdd FILL
XFILL_15_MUX2X1_38 gnd vdd FILL
XFILL_6_AOI21X1_3 gnd vdd FILL
XFILL_15_MUX2X1_49 gnd vdd FILL
XFILL_45_DFFSR_160 gnd vdd FILL
XFILL_22_MUX2X1_5 gnd vdd FILL
XFILL_45_DFFSR_171 gnd vdd FILL
XFILL_45_DFFSR_182 gnd vdd FILL
XFILL_45_DFFSR_193 gnd vdd FILL
XFILL_19_MUX2X1_15 gnd vdd FILL
XFILL_19_MUX2X1_26 gnd vdd FILL
XFILL_19_MUX2X1_37 gnd vdd FILL
XFILL_19_MUX2X1_48 gnd vdd FILL
XFILL_47_DFFSR_2 gnd vdd FILL
XFILL_19_MUX2X1_59 gnd vdd FILL
XNOR3X1_11 NOR3X1_11/A NOR3X1_11/B NOR3X1_11/C gnd NOR3X1_11/Y vdd NOR3X1
XFILL_6_NOR2X1_8 gnd vdd FILL
XFILL_8_MUX2X1_150 gnd vdd FILL
XFILL_8_MUX2X1_161 gnd vdd FILL
XNOR3X1_22 INVX1_26/Y NOR3X1_4/B NOR3X1_6/C gnd NOR3X1_24/B vdd NOR3X1
XNOR3X1_33 NOR3X1_33/A NOR3X1_46/B NOR3X1_46/C gnd NOR3X1_35/A vdd NOR3X1
XFILL_8_MUX2X1_172 gnd vdd FILL
XFILL_7_NOR3X1_19 gnd vdd FILL
XFILL_49_DFFSR_170 gnd vdd FILL
XNOR3X1_44 NOR3X1_44/A NOR3X1_44/B NOR3X1_44/C gnd NOR3X1_44/Y vdd NOR3X1
XFILL_8_MUX2X1_183 gnd vdd FILL
XFILL_49_DFFSR_181 gnd vdd FILL
XFILL_8_MUX2X1_194 gnd vdd FILL
XFILL_49_DFFSR_192 gnd vdd FILL
XFILL_23_DFFSR_106 gnd vdd FILL
XFILL_23_DFFSR_117 gnd vdd FILL
XFILL_23_DFFSR_128 gnd vdd FILL
XFILL_23_DFFSR_139 gnd vdd FILL
XFILL_25_3_1 gnd vdd FILL
XFILL_0_3_1 gnd vdd FILL
XFILL_5_MUX2X1_6 gnd vdd FILL
XFILL_27_DFFSR_105 gnd vdd FILL
XFILL_27_DFFSR_116 gnd vdd FILL
XFILL_27_DFFSR_127 gnd vdd FILL
XFILL_27_DFFSR_138 gnd vdd FILL
XFILL_31_DFFSR_8 gnd vdd FILL
XFILL_27_DFFSR_149 gnd vdd FILL
XFILL_10_NAND3X1_14 gnd vdd FILL
XFILL_10_NAND3X1_25 gnd vdd FILL
XFILL_10_NAND3X1_36 gnd vdd FILL
XFILL_10_NAND3X1_47 gnd vdd FILL
XFILL_10_NAND3X1_58 gnd vdd FILL
XFILL_69_DFFSR_6 gnd vdd FILL
XFILL_10_NAND3X1_69 gnd vdd FILL
XFILL_30_CLKBUF1_14 gnd vdd FILL
XFILL_30_CLKBUF1_25 gnd vdd FILL
XFILL_30_CLKBUF1_36 gnd vdd FILL
XFILL_39_DFFSR_40 gnd vdd FILL
XFILL_39_DFFSR_51 gnd vdd FILL
XFILL_39_DFFSR_62 gnd vdd FILL
XFILL_39_DFFSR_73 gnd vdd FILL
XFILL_39_DFFSR_84 gnd vdd FILL
XFILL_23_NOR3X1_17 gnd vdd FILL
XFILL_39_DFFSR_95 gnd vdd FILL
XFILL_23_NOR3X1_28 gnd vdd FILL
XFILL_23_NOR3X1_39 gnd vdd FILL
XFILL_73_DFFSR_206 gnd vdd FILL
XFILL_73_DFFSR_217 gnd vdd FILL
XFILL_0_DFFSR_14 gnd vdd FILL
XFILL_79_DFFSR_50 gnd vdd FILL
XFILL_73_DFFSR_228 gnd vdd FILL
XFILL_0_DFFSR_25 gnd vdd FILL
XFILL_79_DFFSR_61 gnd vdd FILL
XFILL_0_DFFSR_36 gnd vdd FILL
XFILL_10_NOR2X1_2 gnd vdd FILL
XFILL_73_DFFSR_239 gnd vdd FILL
XFILL_79_DFFSR_72 gnd vdd FILL
XFILL_0_DFFSR_47 gnd vdd FILL
XFILL_79_DFFSR_83 gnd vdd FILL
XFILL_27_NOR3X1_16 gnd vdd FILL
XFILL_27_NOR3X1_27 gnd vdd FILL
XFILL_0_DFFSR_58 gnd vdd FILL
XFILL_79_DFFSR_94 gnd vdd FILL
XFILL_0_DFFSR_69 gnd vdd FILL
XFILL_9_BUFX4_1 gnd vdd FILL
XFILL_27_NOR3X1_38 gnd vdd FILL
XFILL_27_NOR3X1_49 gnd vdd FILL
XFILL_77_DFFSR_205 gnd vdd FILL
XFILL_8_4_1 gnd vdd FILL
XFILL_77_DFFSR_216 gnd vdd FILL
XFILL_77_DFFSR_227 gnd vdd FILL
XFILL_77_DFFSR_238 gnd vdd FILL
XFILL_2_INVX1_90 gnd vdd FILL
XFILL_12_DFFSR_160 gnd vdd FILL
XFILL_19_NOR3X1_2 gnd vdd FILL
XFILL_77_DFFSR_249 gnd vdd FILL
XFILL_2_BUFX2_10 gnd vdd FILL
XFILL_1_CLKBUF1_3 gnd vdd FILL
XFILL_12_DFFSR_171 gnd vdd FILL
XFILL_12_DFFSR_182 gnd vdd FILL
XFILL_12_DFFSR_193 gnd vdd FILL
XFILL_48_DFFSR_60 gnd vdd FILL
XFILL_48_DFFSR_71 gnd vdd FILL
XFILL_48_DFFSR_82 gnd vdd FILL
XFILL_0_NAND3X1_20 gnd vdd FILL
XFILL_48_DFFSR_93 gnd vdd FILL
XFILL_0_NAND3X1_31 gnd vdd FILL
XFILL_0_NAND3X1_42 gnd vdd FILL
XFILL_4_NAND2X1_11 gnd vdd FILL
XFILL_0_NAND3X1_53 gnd vdd FILL
XFILL_16_DFFSR_170 gnd vdd FILL
XFILL_0_NAND3X1_64 gnd vdd FILL
XFILL_4_NAND2X1_22 gnd vdd FILL
XFILL_5_CLKBUF1_2 gnd vdd FILL
XFILL_0_NAND3X1_75 gnd vdd FILL
XFILL_16_DFFSR_181 gnd vdd FILL
XFILL_0_NAND3X1_86 gnd vdd FILL
XFILL_16_DFFSR_192 gnd vdd FILL
XFILL_4_NAND2X1_33 gnd vdd FILL
XFILL_4_NAND2X1_44 gnd vdd FILL
XFILL_0_NAND3X1_97 gnd vdd FILL
XFILL_16_3_1 gnd vdd FILL
XFILL_4_NAND2X1_55 gnd vdd FILL
XFILL_4_NAND2X1_66 gnd vdd FILL
XFILL_4_NAND2X1_77 gnd vdd FILL
XFILL_17_DFFSR_70 gnd vdd FILL
XFILL_4_NAND2X1_88 gnd vdd FILL
XFILL_17_DFFSR_81 gnd vdd FILL
XFILL_17_DFFSR_92 gnd vdd FILL
XFILL_9_CLKBUF1_1 gnd vdd FILL
XFILL_12_CLKBUF1_19 gnd vdd FILL
XFILL_57_DFFSR_80 gnd vdd FILL
XFILL_57_DFFSR_91 gnd vdd FILL
XFILL_62_DFFSR_260 gnd vdd FILL
XFILL_62_DFFSR_271 gnd vdd FILL
XFILL_2_NOR2X1_1 gnd vdd FILL
XFILL_10_NOR2X1_104 gnd vdd FILL
XFILL_9_INVX4_1 gnd vdd FILL
XFILL_10_NOR2X1_115 gnd vdd FILL
XFILL_10_NOR2X1_126 gnd vdd FILL
XFILL_10_NOR2X1_137 gnd vdd FILL
XFILL_66_DFFSR_270 gnd vdd FILL
XFILL_10_NOR2X1_148 gnd vdd FILL
XFILL_10_NOR2X1_159 gnd vdd FILL
XFILL_40_DFFSR_206 gnd vdd FILL
XFILL_26_DFFSR_90 gnd vdd FILL
XFILL_8_AOI21X1_11 gnd vdd FILL
XFILL_40_DFFSR_217 gnd vdd FILL
XFILL_2_OAI21X1_7 gnd vdd FILL
XFILL_8_AOI21X1_22 gnd vdd FILL
XFILL_40_DFFSR_228 gnd vdd FILL
XFILL_8_AOI21X1_33 gnd vdd FILL
XFILL_40_DFFSR_239 gnd vdd FILL
XFILL_8_AOI21X1_44 gnd vdd FILL
XFILL_8_AOI21X1_55 gnd vdd FILL
XFILL_8_AOI21X1_66 gnd vdd FILL
XFILL_18_OAI22X1_13 gnd vdd FILL
XFILL_8_AOI21X1_77 gnd vdd FILL
XFILL_18_OAI22X1_24 gnd vdd FILL
XFILL_18_OAI22X1_35 gnd vdd FILL
XFILL_44_DFFSR_205 gnd vdd FILL
XFILL_18_OAI22X1_46 gnd vdd FILL
XFILL_44_DFFSR_216 gnd vdd FILL
XFILL_3_NOR2X1_20 gnd vdd FILL
XFILL_6_OAI21X1_6 gnd vdd FILL
XFILL_3_NOR2X1_31 gnd vdd FILL
XFILL_3_NOR2X1_42 gnd vdd FILL
XFILL_44_DFFSR_227 gnd vdd FILL
XFILL_66_2_1 gnd vdd FILL
XFILL_3_NOR2X1_53 gnd vdd FILL
XFILL_44_DFFSR_238 gnd vdd FILL
XFILL_44_DFFSR_249 gnd vdd FILL
XFILL_3_NOR2X1_64 gnd vdd FILL
XFILL_2_CLKBUF1_14 gnd vdd FILL
XFILL_2_CLKBUF1_25 gnd vdd FILL
XFILL_3_NOR2X1_75 gnd vdd FILL
XFILL_13_BUFX4_19 gnd vdd FILL
XFILL_3_NOR2X1_86 gnd vdd FILL
XFILL_2_CLKBUF1_36 gnd vdd FILL
XFILL_3_NOR2X1_97 gnd vdd FILL
XFILL_71_DFFSR_105 gnd vdd FILL
XFILL_48_DFFSR_204 gnd vdd FILL
XFILL_9_DFFSR_80 gnd vdd FILL
XFILL_48_DFFSR_215 gnd vdd FILL
XFILL_71_DFFSR_116 gnd vdd FILL
XFILL_7_NOR2X1_30 gnd vdd FILL
XFILL_9_DFFSR_91 gnd vdd FILL
XFILL_71_DFFSR_127 gnd vdd FILL
XFILL_48_DFFSR_226 gnd vdd FILL
XFILL_71_DFFSR_138 gnd vdd FILL
XFILL_7_NOR2X1_41 gnd vdd FILL
XFILL_71_DFFSR_149 gnd vdd FILL
XFILL_7_NOR2X1_52 gnd vdd FILL
XFILL_11_OAI22X1_3 gnd vdd FILL
XFILL_48_DFFSR_237 gnd vdd FILL
XFILL_48_DFFSR_248 gnd vdd FILL
XFILL_7_NOR2X1_63 gnd vdd FILL
XFILL_48_DFFSR_259 gnd vdd FILL
XFILL_7_NOR2X1_74 gnd vdd FILL
XFILL_7_NOR2X1_85 gnd vdd FILL
XFILL_75_DFFSR_104 gnd vdd FILL
XFILL_7_NOR2X1_96 gnd vdd FILL
XFILL_0_NOR2X1_110 gnd vdd FILL
XFILL_11_OAI21X1_15 gnd vdd FILL
XFILL_75_DFFSR_115 gnd vdd FILL
XFILL_50_6_2 gnd vdd FILL
XFILL_11_OAI21X1_26 gnd vdd FILL
XFILL_75_DFFSR_126 gnd vdd FILL
XFILL_0_NOR2X1_121 gnd vdd FILL
XFILL_75_DFFSR_137 gnd vdd FILL
XFILL_0_NOR2X1_132 gnd vdd FILL
XFILL_0_DFFSR_7 gnd vdd FILL
XFILL_15_OAI22X1_2 gnd vdd FILL
XFILL_75_DFFSR_148 gnd vdd FILL
XFILL_0_NOR2X1_143 gnd vdd FILL
XFILL_11_OAI21X1_37 gnd vdd FILL
XFILL_11_OAI21X1_48 gnd vdd FILL
XFILL_0_NOR2X1_154 gnd vdd FILL
XFILL_13_DFFSR_5 gnd vdd FILL
XFILL_75_DFFSR_159 gnd vdd FILL
XFILL_0_NOR2X1_165 gnd vdd FILL
XFILL_0_NOR2X1_176 gnd vdd FILL
XFILL_70_DFFSR_6 gnd vdd FILL
XFILL_0_NOR2X1_187 gnd vdd FILL
XFILL_79_DFFSR_103 gnd vdd FILL
XFILL_0_NOR2X1_198 gnd vdd FILL
XFILL_79_DFFSR_114 gnd vdd FILL
XFILL_79_DFFSR_125 gnd vdd FILL
XFILL_79_DFFSR_136 gnd vdd FILL
XFILL_19_OAI22X1_1 gnd vdd FILL
XFILL_79_DFFSR_147 gnd vdd FILL
XFILL_79_DFFSR_158 gnd vdd FILL
XFILL_10_NAND2X1_80 gnd vdd FILL
XFILL_8_OAI22X1_30 gnd vdd FILL
XFILL_10_NAND2X1_91 gnd vdd FILL
XFILL_79_DFFSR_169 gnd vdd FILL
XFILL_8_OAI22X1_41 gnd vdd FILL
XBUFX2_4 INVX2_4/A gnd addr[0] vdd BUFX2
XFILL_33_DFFSR_270 gnd vdd FILL
XFILL_0_MUX2X1_105 gnd vdd FILL
XFILL_0_MUX2X1_116 gnd vdd FILL
XFILL_3_NAND2X1_8 gnd vdd FILL
XFILL_0_MUX2X1_127 gnd vdd FILL
XFILL_0_MUX2X1_138 gnd vdd FILL
XFILL_35_DFFSR_9 gnd vdd FILL
XFILL_0_MUX2X1_149 gnd vdd FILL
XFILL_5_BUFX4_18 gnd vdd FILL
XFILL_5_BUFX4_29 gnd vdd FILL
XFILL_58_7_2 gnd vdd FILL
XFILL_60_DFFSR_170 gnd vdd FILL
XFILL_1_OAI21X1_10 gnd vdd FILL
XFILL_60_DFFSR_181 gnd vdd FILL
XFILL_1_OAI21X1_21 gnd vdd FILL
XFILL_60_DFFSR_192 gnd vdd FILL
XFILL_7_NAND2X1_7 gnd vdd FILL
XFILL_57_2_1 gnd vdd FILL
XFILL_11_DFFSR_205 gnd vdd FILL
XFILL_1_OAI21X1_32 gnd vdd FILL
XFILL_1_OAI21X1_43 gnd vdd FILL
XFILL_11_DFFSR_216 gnd vdd FILL
XFILL_3_MUX2X1_60 gnd vdd FILL
XFILL_11_DFFSR_227 gnd vdd FILL
XFILL_3_MUX2X1_71 gnd vdd FILL
XFILL_11_DFFSR_238 gnd vdd FILL
XFILL_11_DFFSR_249 gnd vdd FILL
XFILL_3_MUX2X1_82 gnd vdd FILL
XFILL_3_MUX2X1_93 gnd vdd FILL
XFILL_64_DFFSR_180 gnd vdd FILL
XFILL_64_DFFSR_191 gnd vdd FILL
XFILL_15_DFFSR_204 gnd vdd FILL
XFILL_15_DFFSR_215 gnd vdd FILL
XFILL_12_NAND3X1_4 gnd vdd FILL
XFILL_14_AOI21X1_80 gnd vdd FILL
XFILL_7_MUX2X1_70 gnd vdd FILL
XFILL_15_DFFSR_226 gnd vdd FILL
XFILL_15_DFFSR_237 gnd vdd FILL
XFILL_7_MUX2X1_81 gnd vdd FILL
XFILL_15_DFFSR_248 gnd vdd FILL
XFILL_7_MUX2X1_92 gnd vdd FILL
XFILL_15_DFFSR_259 gnd vdd FILL
XFILL_41_6_2 gnd vdd FILL
XFILL_68_DFFSR_190 gnd vdd FILL
XFILL_42_DFFSR_104 gnd vdd FILL
XFILL_40_1_1 gnd vdd FILL
XFILL_19_DFFSR_203 gnd vdd FILL
XFILL_12_AND2X2_6 gnd vdd FILL
XFILL_42_DFFSR_115 gnd vdd FILL
XFILL_19_DFFSR_214 gnd vdd FILL
XFILL_42_DFFSR_126 gnd vdd FILL
XFILL_19_DFFSR_225 gnd vdd FILL
XFILL_42_DFFSR_137 gnd vdd FILL
XINVX2_4 INVX2_4/A gnd INVX2_4/Y vdd INVX2
XFILL_42_DFFSR_148 gnd vdd FILL
XFILL_19_DFFSR_236 gnd vdd FILL
XFILL_19_DFFSR_247 gnd vdd FILL
XFILL_19_DFFSR_258 gnd vdd FILL
XFILL_42_DFFSR_159 gnd vdd FILL
XFILL_19_DFFSR_269 gnd vdd FILL
XFILL_46_DFFSR_103 gnd vdd FILL
XFILL_46_DFFSR_114 gnd vdd FILL
XAOI21X1_4 BUFX4_80/Y AOI21X1_7/B AOI21X1_4/C gnd DFFSR_139/D vdd AOI21X1
XFILL_3_NAND3X1_19 gnd vdd FILL
XFILL_46_DFFSR_125 gnd vdd FILL
XFILL_46_DFFSR_136 gnd vdd FILL
XFILL_46_DFFSR_147 gnd vdd FILL
XFILL_46_DFFSR_158 gnd vdd FILL
XFILL_46_DFFSR_169 gnd vdd FILL
XMUX2X1_140 BUFX4_66/Y NOR3X1_14/A AOI21X1_1/B gnd DFFSR_180/D vdd MUX2X1
XMUX2X1_151 BUFX4_93/Y NOR3X1_41/A AOI21X1_1/B gnd DFFSR_182/D vdd MUX2X1
XMUX2X1_162 BUFX4_81/Y OAI22X1_4/C MUX2X1_2/S gnd DFFSR_174/D vdd MUX2X1
XMUX2X1_173 BUFX4_68/Y INVX1_13/Y MUX2X1_2/S gnd DFFSR_175/D vdd MUX2X1
XFILL_17_MUX2X1_130 gnd vdd FILL
XFILL_12_AOI22X1_9 gnd vdd FILL
XFILL_17_MUX2X1_141 gnd vdd FILL
XMUX2X1_184 BUFX4_78/Y INVX1_24/Y MUX2X1_2/S gnd DFFSR_176/D vdd MUX2X1
XFILL_17_MUX2X1_152 gnd vdd FILL
XFILL_17_MUX2X1_163 gnd vdd FILL
XFILL_23_MUX2X1_90 gnd vdd FILL
XFILL_17_MUX2X1_174 gnd vdd FILL
XFILL_17_MUX2X1_185 gnd vdd FILL
XFILL_49_7_2 gnd vdd FILL
XFILL_16_AOI22X1_8 gnd vdd FILL
XFILL_48_2_1 gnd vdd FILL
XINVX1_80 INVX1_80/A gnd INVX1_80/Y vdd INVX1
XINVX1_91 INVX1_91/A gnd INVX1_91/Y vdd INVX1
XFILL_54_8 gnd vdd FILL
XFILL_3_INVX1_13 gnd vdd FILL
XFILL_3_INVX1_24 gnd vdd FILL
XFILL_10_INVX8_3 gnd vdd FILL
XFILL_3_INVX1_35 gnd vdd FILL
XFILL_3_INVX1_46 gnd vdd FILL
XFILL_4_AND2X2_5 gnd vdd FILL
XFILL_3_INVX1_57 gnd vdd FILL
XFILL_31_DFFSR_180 gnd vdd FILL
XFILL_3_INVX1_68 gnd vdd FILL
XFILL_49_DFFSR_16 gnd vdd FILL
XFILL_31_DFFSR_191 gnd vdd FILL
XFILL_3_INVX1_79 gnd vdd FILL
XFILL_49_DFFSR_27 gnd vdd FILL
XFILL_49_DFFSR_38 gnd vdd FILL
XFILL_49_DFFSR_49 gnd vdd FILL
XFILL_32_6_2 gnd vdd FILL
XFILL_31_1_1 gnd vdd FILL
XFILL_35_DFFSR_190 gnd vdd FILL
XFILL_1_BUFX4_11 gnd vdd FILL
XFILL_52_DFFSR_3 gnd vdd FILL
XFILL_1_BUFX4_22 gnd vdd FILL
XFILL_1_BUFX4_33 gnd vdd FILL
XFILL_1_BUFX4_44 gnd vdd FILL
XFILL_18_DFFSR_15 gnd vdd FILL
XFILL_18_DFFSR_26 gnd vdd FILL
XFILL_1_BUFX4_55 gnd vdd FILL
XFILL_1_BUFX4_66 gnd vdd FILL
XFILL_18_DFFSR_37 gnd vdd FILL
XFILL_7_MUX2X1_180 gnd vdd FILL
XFILL_1_BUFX4_77 gnd vdd FILL
XFILL_18_DFFSR_48 gnd vdd FILL
XFILL_1_BUFX4_88 gnd vdd FILL
XFILL_13_DFFSR_103 gnd vdd FILL
XFILL_18_DFFSR_59 gnd vdd FILL
XFILL_7_MUX2X1_191 gnd vdd FILL
XFILL_1_BUFX4_99 gnd vdd FILL
XFILL_13_DFFSR_114 gnd vdd FILL
XFILL_13_DFFSR_125 gnd vdd FILL
XFILL_13_DFFSR_136 gnd vdd FILL
XFILL_58_DFFSR_14 gnd vdd FILL
XFILL_13_DFFSR_147 gnd vdd FILL
XNOR2X1_2 NOR2X1_2/A NOR2X1_2/B gnd NOR2X1_2/Y vdd NOR2X1
XFILL_58_DFFSR_25 gnd vdd FILL
XFILL_13_DFFSR_158 gnd vdd FILL
XFILL_58_DFFSR_36 gnd vdd FILL
XFILL_13_DFFSR_169 gnd vdd FILL
XFILL_58_DFFSR_47 gnd vdd FILL
XFILL_17_DFFSR_102 gnd vdd FILL
XFILL_58_DFFSR_58 gnd vdd FILL
XFILL_58_DFFSR_69 gnd vdd FILL
XFILL_3_NOR2X1_109 gnd vdd FILL
XFILL_17_DFFSR_113 gnd vdd FILL
XFILL_17_DFFSR_124 gnd vdd FILL
XFILL_17_DFFSR_135 gnd vdd FILL
XFILL_17_DFFSR_146 gnd vdd FILL
XFILL_4_DFFSR_8 gnd vdd FILL
XFILL_17_DFFSR_157 gnd vdd FILL
XFILL_17_DFFSR_6 gnd vdd FILL
XFILL_17_DFFSR_168 gnd vdd FILL
XFILL_17_DFFSR_179 gnd vdd FILL
XFILL_74_DFFSR_7 gnd vdd FILL
XFILL_27_DFFSR_13 gnd vdd FILL
XFILL_27_DFFSR_24 gnd vdd FILL
XFILL_27_DFFSR_35 gnd vdd FILL
XFILL_39_2_1 gnd vdd FILL
XFILL_27_DFFSR_46 gnd vdd FILL
XFILL_27_DFFSR_57 gnd vdd FILL
XFILL_27_DFFSR_68 gnd vdd FILL
XFILL_27_DFFSR_79 gnd vdd FILL
XFILL_13_NOR3X1_14 gnd vdd FILL
XFILL_67_DFFSR_12 gnd vdd FILL
XFILL_13_NOR3X1_25 gnd vdd FILL
XFILL_67_DFFSR_23 gnd vdd FILL
XFILL_13_NOR3X1_36 gnd vdd FILL
XFILL_67_DFFSR_34 gnd vdd FILL
XFILL_13_NOR3X1_47 gnd vdd FILL
XFILL_63_DFFSR_203 gnd vdd FILL
XFILL_67_DFFSR_45 gnd vdd FILL
XFILL_67_DFFSR_56 gnd vdd FILL
XFILL_63_DFFSR_214 gnd vdd FILL
XFILL_63_DFFSR_225 gnd vdd FILL
XFILL_67_DFFSR_67 gnd vdd FILL
XFILL_6_BUFX4_105 gnd vdd FILL
XFILL_67_DFFSR_78 gnd vdd FILL
XFILL_63_DFFSR_236 gnd vdd FILL
XFILL_67_DFFSR_89 gnd vdd FILL
XFILL_63_DFFSR_247 gnd vdd FILL
XFILL_17_NOR3X1_13 gnd vdd FILL
XFILL_63_DFFSR_258 gnd vdd FILL
XFILL_63_DFFSR_269 gnd vdd FILL
XFILL_17_NOR3X1_24 gnd vdd FILL
XFILL_23_6_2 gnd vdd FILL
XFILL_17_NOR3X1_35 gnd vdd FILL
XFILL_67_DFFSR_202 gnd vdd FILL
XFILL_17_NOR3X1_46 gnd vdd FILL
XFILL_22_1_1 gnd vdd FILL
XFILL_67_DFFSR_213 gnd vdd FILL
XFILL_36_DFFSR_11 gnd vdd FILL
XFILL_67_DFFSR_224 gnd vdd FILL
XFILL_0_OAI22X1_18 gnd vdd FILL
XFILL_36_DFFSR_22 gnd vdd FILL
XFILL_67_DFFSR_235 gnd vdd FILL
XFILL_36_DFFSR_33 gnd vdd FILL
XFILL_0_OAI22X1_29 gnd vdd FILL
XFILL_67_DFFSR_246 gnd vdd FILL
XFILL_36_DFFSR_44 gnd vdd FILL
XFILL_36_DFFSR_55 gnd vdd FILL
XFILL_67_DFFSR_257 gnd vdd FILL
XFILL_67_DFFSR_268 gnd vdd FILL
XFILL_36_DFFSR_66 gnd vdd FILL
XFILL_22_CLKBUF1_9 gnd vdd FILL
XFILL_36_DFFSR_77 gnd vdd FILL
XAOI21X1_12 BUFX4_72/Y NOR2X1_2/B NOR2X1_2/Y gnd DFFSR_172/D vdd AOI21X1
XFILL_13_AOI22X1_11 gnd vdd FILL
XFILL_36_DFFSR_88 gnd vdd FILL
XFILL_0_NOR2X1_19 gnd vdd FILL
XFILL_36_DFFSR_99 gnd vdd FILL
XFILL_76_DFFSR_10 gnd vdd FILL
XAOI21X1_23 BUFX4_72/Y NOR2X1_46/B NOR2X1_46/Y gnd DFFSR_167/D vdd AOI21X1
XAOI21X1_34 BUFX4_81/Y NOR2X1_90/B NOR2X1_79/Y gnd DFFSR_156/D vdd AOI21X1
XFILL_76_DFFSR_21 gnd vdd FILL
XAOI21X1_45 MUX2X1_1/A NOR2X1_90/B NOR2X1_90/Y gnd DFFSR_158/D vdd AOI21X1
XAOI21X1_56 BUFX4_76/Y NOR2X1_90/B NOR2X1_101/Y gnd DFFSR_159/D vdd AOI21X1
XFILL_76_DFFSR_32 gnd vdd FILL
XAOI21X1_67 MUX2X1_2/A NOR2X1_90/B NOR2X1_113/Y gnd DFFSR_160/D vdd AOI21X1
XFILL_76_DFFSR_43 gnd vdd FILL
XFILL_76_DFFSR_54 gnd vdd FILL
XAOI21X1_78 BUFX4_83/Y AOI21X1_3/B NOR2X1_124/Y gnd DFFSR_148/D vdd AOI21X1
XFILL_76_DFFSR_65 gnd vdd FILL
XFILL_3_NAND2X1_30 gnd vdd FILL
XFILL_76_DFFSR_76 gnd vdd FILL
XFILL_26_CLKBUF1_8 gnd vdd FILL
XFILL_3_NAND2X1_41 gnd vdd FILL
XFILL_3_NAND2X1_52 gnd vdd FILL
XFILL_76_DFFSR_87 gnd vdd FILL
XFILL_4_NOR2X1_18 gnd vdd FILL
XFILL_76_DFFSR_98 gnd vdd FILL
XOAI21X1_7 OAI21X1_7/A OAI21X1_7/B OAI21X1_7/C gnd OAI21X1_7/Y vdd OAI21X1
XFILL_3_NAND2X1_63 gnd vdd FILL
XFILL_3_NAND2X1_74 gnd vdd FILL
XFILL_4_NOR2X1_29 gnd vdd FILL
XFILL_11_BUFX4_6 gnd vdd FILL
XFILL_3_NAND2X1_85 gnd vdd FILL
XFILL_3_NAND2X1_96 gnd vdd FILL
XFILL_45_DFFSR_20 gnd vdd FILL
XFILL_45_DFFSR_31 gnd vdd FILL
XFILL_16_NOR3X1_6 gnd vdd FILL
XFILL_11_CLKBUF1_16 gnd vdd FILL
XFILL_45_DFFSR_42 gnd vdd FILL
XFILL_8_NOR2X1_17 gnd vdd FILL
XFILL_45_DFFSR_53 gnd vdd FILL
XFILL_11_CLKBUF1_27 gnd vdd FILL
XFILL_11_CLKBUF1_38 gnd vdd FILL
XFILL_8_NOR2X1_28 gnd vdd FILL
XFILL_45_DFFSR_64 gnd vdd FILL
XFILL_45_DFFSR_75 gnd vdd FILL
XFILL_8_NOR2X1_39 gnd vdd FILL
XFILL_45_DFFSR_86 gnd vdd FILL
XFILL_6_7_2 gnd vdd FILL
XFILL_5_2_1 gnd vdd FILL
XFILL_45_DFFSR_97 gnd vdd FILL
XFILL_85_DFFSR_30 gnd vdd FILL
XFILL_85_DFFSR_41 gnd vdd FILL
XFILL_85_DFFSR_52 gnd vdd FILL
XFILL_85_DFFSR_63 gnd vdd FILL
XFILL_85_DFFSR_74 gnd vdd FILL
XFILL_14_DFFSR_30 gnd vdd FILL
XFILL_85_DFFSR_85 gnd vdd FILL
XFILL_29_CLKBUF1_40 gnd vdd FILL
XFILL_14_DFFSR_41 gnd vdd FILL
XFILL_85_DFFSR_96 gnd vdd FILL
XFILL_14_DFFSR_52 gnd vdd FILL
XFILL_14_DFFSR_63 gnd vdd FILL
XFILL_14_DFFSR_74 gnd vdd FILL
XFILL_14_DFFSR_85 gnd vdd FILL
XFILL_14_DFFSR_96 gnd vdd FILL
XFILL_30_DFFSR_203 gnd vdd FILL
XFILL_30_DFFSR_214 gnd vdd FILL
XFILL_14_6_2 gnd vdd FILL
XOAI22X1_20 INVX1_42/Y INVX1_121/A INVX1_44/Y INVX1_120/A gnd NOR3X1_30/C vdd OAI22X1
XFILL_7_AOI21X1_30 gnd vdd FILL
XFILL_54_DFFSR_40 gnd vdd FILL
XFILL_30_DFFSR_225 gnd vdd FILL
XFILL_25_NOR3X1_4 gnd vdd FILL
XFILL_54_DFFSR_51 gnd vdd FILL
XOAI22X1_31 INVX1_5/Y OAI22X1_5/B INVX1_10/Y OAI22X1_5/D gnd NOR2X1_94/B vdd OAI22X1
XFILL_30_DFFSR_236 gnd vdd FILL
XOAI22X1_42 INVX1_92/Y OAI22X1_6/B INVX1_95/Y OAI22X1_6/D gnd OAI22X1_42/Y vdd OAI22X1
XFILL_7_AOI21X1_41 gnd vdd FILL
XFILL_30_DFFSR_247 gnd vdd FILL
XFILL_13_1_1 gnd vdd FILL
XFILL_7_AOI21X1_52 gnd vdd FILL
XFILL_30_DFFSR_258 gnd vdd FILL
XFILL_54_DFFSR_62 gnd vdd FILL
XFILL_17_OAI22X1_10 gnd vdd FILL
XFILL_30_DFFSR_269 gnd vdd FILL
XFILL_54_DFFSR_73 gnd vdd FILL
XFILL_7_AOI21X1_63 gnd vdd FILL
XFILL_54_DFFSR_84 gnd vdd FILL
XFILL_7_AOI21X1_74 gnd vdd FILL
XFILL_17_OAI22X1_21 gnd vdd FILL
XFILL_54_DFFSR_95 gnd vdd FILL
XFILL_17_OAI22X1_32 gnd vdd FILL
XFILL_34_DFFSR_202 gnd vdd FILL
XFILL_17_OAI22X1_43 gnd vdd FILL
XFILL_34_DFFSR_213 gnd vdd FILL
XFILL_34_DFFSR_224 gnd vdd FILL
XFILL_34_DFFSR_235 gnd vdd FILL
XFILL_34_DFFSR_246 gnd vdd FILL
XFILL_1_CLKBUF1_11 gnd vdd FILL
XFILL_3_DFFSR_270 gnd vdd FILL
XFILL_34_DFFSR_257 gnd vdd FILL
XFILL_1_CLKBUF1_22 gnd vdd FILL
XFILL_34_DFFSR_268 gnd vdd FILL
XFILL_1_CLKBUF1_33 gnd vdd FILL
XFILL_0_MUX2X1_15 gnd vdd FILL
XFILL_61_DFFSR_102 gnd vdd FILL
XFILL_0_MUX2X1_26 gnd vdd FILL
XFILL_23_DFFSR_50 gnd vdd FILL
XFILL_38_DFFSR_201 gnd vdd FILL
XFILL_0_MUX2X1_37 gnd vdd FILL
XFILL_23_DFFSR_61 gnd vdd FILL
XFILL_38_DFFSR_212 gnd vdd FILL
XFILL_0_MUX2X1_48 gnd vdd FILL
XFILL_61_DFFSR_113 gnd vdd FILL
XFILL_61_DFFSR_124 gnd vdd FILL
XFILL_14_INVX8_4 gnd vdd FILL
XFILL_38_DFFSR_223 gnd vdd FILL
XFILL_23_DFFSR_72 gnd vdd FILL
XFILL_23_DFFSR_83 gnd vdd FILL
XFILL_38_DFFSR_234 gnd vdd FILL
XFILL_61_DFFSR_135 gnd vdd FILL
XFILL_0_MUX2X1_59 gnd vdd FILL
XFILL_61_DFFSR_146 gnd vdd FILL
XFILL_23_DFFSR_94 gnd vdd FILL
XFILL_61_DFFSR_157 gnd vdd FILL
XFILL_38_DFFSR_245 gnd vdd FILL
XFILL_8_NOR3X1_5 gnd vdd FILL
XFILL_38_DFFSR_256 gnd vdd FILL
XFILL_38_DFFSR_267 gnd vdd FILL
XFILL_61_DFFSR_168 gnd vdd FILL
XFILL_4_MUX2X1_14 gnd vdd FILL
XFILL_61_DFFSR_179 gnd vdd FILL
XFILL_4_MUX2X1_25 gnd vdd FILL
XFILL_65_DFFSR_101 gnd vdd FILL
XFILL_63_DFFSR_60 gnd vdd FILL
XFILL_4_MUX2X1_36 gnd vdd FILL
XFILL_65_DFFSR_112 gnd vdd FILL
XFILL_4_MUX2X1_47 gnd vdd FILL
XFILL_10_OAI21X1_12 gnd vdd FILL
XFILL_63_DFFSR_71 gnd vdd FILL
XFILL_4_MUX2X1_58 gnd vdd FILL
XFILL_10_OAI21X1_23 gnd vdd FILL
XFILL_65_DFFSR_123 gnd vdd FILL
XFILL_63_DFFSR_82 gnd vdd FILL
XFILL_65_DFFSR_134 gnd vdd FILL
XFILL_10_OAI21X1_34 gnd vdd FILL
XFILL_4_MUX2X1_69 gnd vdd FILL
XFILL_63_DFFSR_93 gnd vdd FILL
XFILL_65_DFFSR_145 gnd vdd FILL
XFILL_65_DFFSR_156 gnd vdd FILL
XFILL_3_4 gnd vdd FILL
XFILL_10_OAI21X1_45 gnd vdd FILL
XFILL_8_MUX2X1_13 gnd vdd FILL
XFILL_65_DFFSR_167 gnd vdd FILL
XFILL_65_DFFSR_178 gnd vdd FILL
XFILL_69_DFFSR_100 gnd vdd FILL
XFILL_65_DFFSR_189 gnd vdd FILL
XFILL_8_MUX2X1_24 gnd vdd FILL
XFILL_56_DFFSR_4 gnd vdd FILL
XFILL_6_DFFSR_40 gnd vdd FILL
XFILL_8_MUX2X1_35 gnd vdd FILL
XFILL_69_DFFSR_111 gnd vdd FILL
XFILL_6_DFFSR_51 gnd vdd FILL
XFILL_69_DFFSR_122 gnd vdd FILL
XFILL_8_MUX2X1_46 gnd vdd FILL
XFILL_6_DFFSR_62 gnd vdd FILL
XFILL_8_MUX2X1_57 gnd vdd FILL
XFILL_69_DFFSR_133 gnd vdd FILL
XFILL_8_MUX2X1_68 gnd vdd FILL
XFILL_69_DFFSR_144 gnd vdd FILL
XFILL_6_DFFSR_73 gnd vdd FILL
XFILL_12_OAI21X1_1 gnd vdd FILL
XFILL_8_MUX2X1_79 gnd vdd FILL
XFILL_6_DFFSR_84 gnd vdd FILL
XFILL_69_DFFSR_155 gnd vdd FILL
XFILL_6_DFFSR_95 gnd vdd FILL
XFILL_32_DFFSR_70 gnd vdd FILL
XFILL_69_DFFSR_166 gnd vdd FILL
XFILL_32_DFFSR_81 gnd vdd FILL
XFILL_64_5_2 gnd vdd FILL
XFILL_69_DFFSR_177 gnd vdd FILL
XFILL_32_DFFSR_92 gnd vdd FILL
XFILL_69_DFFSR_188 gnd vdd FILL
XFILL_45_4 gnd vdd FILL
XFILL_69_DFFSR_199 gnd vdd FILL
XFILL_63_0_1 gnd vdd FILL
XFILL_38_3 gnd vdd FILL
XFILL_72_DFFSR_80 gnd vdd FILL
XFILL_72_DFFSR_91 gnd vdd FILL
XFILL_20_MUX2X1_12 gnd vdd FILL
XFILL_20_MUX2X1_23 gnd vdd FILL
XFILL_20_MUX2X1_34 gnd vdd FILL
XFILL_8_DFFSR_9 gnd vdd FILL
XFILL_20_MUX2X1_45 gnd vdd FILL
XFILL_20_MUX2X1_56 gnd vdd FILL
XFILL_20_MUX2X1_67 gnd vdd FILL
XFILL_20_MUX2X1_78 gnd vdd FILL
XFILL_78_DFFSR_8 gnd vdd FILL
XFILL_20_MUX2X1_89 gnd vdd FILL
XFILL_0_OAI21X1_40 gnd vdd FILL
XFILL_41_DFFSR_90 gnd vdd FILL
XFILL_32_DFFSR_101 gnd vdd FILL
XFILL_32_DFFSR_112 gnd vdd FILL
XFILL_32_DFFSR_123 gnd vdd FILL
XFILL_32_DFFSR_134 gnd vdd FILL
XFILL_32_DFFSR_145 gnd vdd FILL
XFILL_32_DFFSR_156 gnd vdd FILL
XFILL_1_DFFSR_180 gnd vdd FILL
XFILL_32_DFFSR_167 gnd vdd FILL
XFILL_32_DFFSR_178 gnd vdd FILL
XFILL_1_DFFSR_191 gnd vdd FILL
XFILL_36_DFFSR_100 gnd vdd FILL
XFILL_32_DFFSR_189 gnd vdd FILL
XFILL_36_DFFSR_111 gnd vdd FILL
XFILL_2_NAND3X1_16 gnd vdd FILL
XFILL_36_DFFSR_122 gnd vdd FILL
XFILL_36_DFFSR_133 gnd vdd FILL
XFILL_2_NAND3X1_27 gnd vdd FILL
XFILL_55_5_2 gnd vdd FILL
XFILL_36_DFFSR_144 gnd vdd FILL
XFILL_2_NAND3X1_38 gnd vdd FILL
XFILL_36_DFFSR_155 gnd vdd FILL
XFILL_2_NAND3X1_49 gnd vdd FILL
XFILL_36_DFFSR_166 gnd vdd FILL
XFILL_54_0_1 gnd vdd FILL
XFILL_6_NAND2X1_18 gnd vdd FILL
XFILL_36_DFFSR_177 gnd vdd FILL
XFILL_5_DFFSR_190 gnd vdd FILL
XFILL_6_NAND2X1_29 gnd vdd FILL
XFILL_36_DFFSR_188 gnd vdd FILL
XFILL_2_BUFX4_9 gnd vdd FILL
XFILL_36_DFFSR_199 gnd vdd FILL
XFILL_15_BUFX4_7 gnd vdd FILL
XFILL_16_MUX2X1_160 gnd vdd FILL
XFILL_16_MUX2X1_171 gnd vdd FILL
XFILL_16_MUX2X1_182 gnd vdd FILL
XFILL_82_DFFSR_201 gnd vdd FILL
XFILL_16_MUX2X1_193 gnd vdd FILL
XFILL_82_DFFSR_212 gnd vdd FILL
XFILL_82_DFFSR_223 gnd vdd FILL
XFILL_82_DFFSR_234 gnd vdd FILL
XFILL_82_DFFSR_245 gnd vdd FILL
XFILL_82_DFFSR_256 gnd vdd FILL
XFILL_82_DFFSR_267 gnd vdd FILL
XFILL_86_DFFSR_200 gnd vdd FILL
XFILL_86_DFFSR_211 gnd vdd FILL
XFILL_86_DFFSR_222 gnd vdd FILL
XFILL_13_AOI21X1_7 gnd vdd FILL
XFILL_86_DFFSR_233 gnd vdd FILL
XFILL_86_DFFSR_244 gnd vdd FILL
XFILL_86_DFFSR_255 gnd vdd FILL
XFILL_86_DFFSR_266 gnd vdd FILL
XFILL_11_BUFX2_3 gnd vdd FILL
XFILL_2_INVX1_150 gnd vdd FILL
XFILL_2_INVX1_161 gnd vdd FILL
XFILL_2_INVX1_172 gnd vdd FILL
XFILL_2_INVX1_183 gnd vdd FILL
XFILL_2_INVX1_194 gnd vdd FILL
XFILL_21_CLKBUF1_17 gnd vdd FILL
XFILL_21_CLKBUF1_28 gnd vdd FILL
XFILL_21_CLKBUF1_39 gnd vdd FILL
XFILL_6_INVX1_160 gnd vdd FILL
XFILL_38_DFFSR_1 gnd vdd FILL
XFILL_6_INVX1_171 gnd vdd FILL
XFILL_0_INVX1_17 gnd vdd FILL
XFILL_6_INVX1_182 gnd vdd FILL
XFILL_0_INVX1_28 gnd vdd FILL
XFILL_6_INVX1_193 gnd vdd FILL
XFILL_0_INVX1_39 gnd vdd FILL
XFILL_46_5_2 gnd vdd FILL
XFILL_45_0_1 gnd vdd FILL
XFILL_0_OAI22X1_1 gnd vdd FILL
XFILL_2_NOR2X1_106 gnd vdd FILL
XFILL_24_9 gnd vdd FILL
XFILL_2_NOR2X1_117 gnd vdd FILL
XFILL_86_DFFSR_19 gnd vdd FILL
XFILL_2_NOR2X1_128 gnd vdd FILL
XFILL_2_NOR2X1_139 gnd vdd FILL
XFILL_22_DFFSR_7 gnd vdd FILL
XFILL_15_DFFSR_19 gnd vdd FILL
XFILL_55_DFFSR_18 gnd vdd FILL
XFILL_55_DFFSR_29 gnd vdd FILL
XFILL_53_DFFSR_200 gnd vdd FILL
XFILL_53_DFFSR_211 gnd vdd FILL
XFILL_53_DFFSR_222 gnd vdd FILL
XFILL_53_DFFSR_233 gnd vdd FILL
XFILL_53_DFFSR_244 gnd vdd FILL
XFILL_53_DFFSR_255 gnd vdd FILL
XFILL_53_DFFSR_266 gnd vdd FILL
XFILL_80_DFFSR_100 gnd vdd FILL
XFILL_9_NAND3X1_80 gnd vdd FILL
XFILL_9_NAND3X1_91 gnd vdd FILL
XFILL_57_DFFSR_210 gnd vdd FILL
XFILL_24_DFFSR_17 gnd vdd FILL
XFILL_80_DFFSR_111 gnd vdd FILL
XFILL_7_NOR2X1_206 gnd vdd FILL
XFILL_24_DFFSR_28 gnd vdd FILL
XFILL_1_1 gnd vdd FILL
XFILL_57_DFFSR_221 gnd vdd FILL
XFILL_80_DFFSR_122 gnd vdd FILL
XFILL_80_DFFSR_133 gnd vdd FILL
XFILL_15_BUFX4_60 gnd vdd FILL
XFILL_24_DFFSR_39 gnd vdd FILL
XFILL_57_DFFSR_232 gnd vdd FILL
XFILL_80_DFFSR_144 gnd vdd FILL
XFILL_15_BUFX4_71 gnd vdd FILL
XFILL_57_DFFSR_243 gnd vdd FILL
XFILL_80_DFFSR_155 gnd vdd FILL
XFILL_15_BUFX4_82 gnd vdd FILL
XFILL_57_DFFSR_254 gnd vdd FILL
XFILL_15_BUFX4_93 gnd vdd FILL
XFILL_80_DFFSR_166 gnd vdd FILL
XFILL_57_DFFSR_265 gnd vdd FILL
XFILL_80_DFFSR_177 gnd vdd FILL
XFILL_12_CLKBUF1_6 gnd vdd FILL
XFILL_3_OAI21X1_17 gnd vdd FILL
XFILL_80_DFFSR_188 gnd vdd FILL
XFILL_0_DFFSR_203 gnd vdd FILL
XFILL_3_OAI21X1_28 gnd vdd FILL
XFILL_84_DFFSR_110 gnd vdd FILL
XFILL_80_DFFSR_199 gnd vdd FILL
XFILL_0_DFFSR_214 gnd vdd FILL
XFILL_64_DFFSR_16 gnd vdd FILL
XFILL_3_OAI21X1_39 gnd vdd FILL
XFILL_0_DFFSR_225 gnd vdd FILL
XFILL_50_2 gnd vdd FILL
XFILL_64_DFFSR_27 gnd vdd FILL
XFILL_84_DFFSR_121 gnd vdd FILL
XFILL_84_DFFSR_132 gnd vdd FILL
XFILL_37_5_2 gnd vdd FILL
XFILL_64_DFFSR_38 gnd vdd FILL
XFILL_0_DFFSR_236 gnd vdd FILL
XFILL_84_DFFSR_143 gnd vdd FILL
XFILL_0_DFFSR_247 gnd vdd FILL
XFILL_64_DFFSR_49 gnd vdd FILL
XFILL_84_DFFSR_154 gnd vdd FILL
XFILL_0_DFFSR_258 gnd vdd FILL
XFILL_0_DFFSR_269 gnd vdd FILL
XFILL_36_0_1 gnd vdd FILL
XFILL_84_DFFSR_165 gnd vdd FILL
XFILL_43_1 gnd vdd FILL
XFILL_84_DFFSR_176 gnd vdd FILL
XFILL_16_CLKBUF1_5 gnd vdd FILL
XFILL_4_DFFSR_202 gnd vdd FILL
XFILL_84_DFFSR_187 gnd vdd FILL
XFILL_4_DFFSR_213 gnd vdd FILL
XFILL_84_DFFSR_198 gnd vdd FILL
XFILL_1_NAND3X1_2 gnd vdd FILL
XFILL_2_NAND2X1_60 gnd vdd FILL
XFILL_4_DFFSR_224 gnd vdd FILL
XFILL_2_NAND2X1_71 gnd vdd FILL
XFILL_4_DFFSR_235 gnd vdd FILL
XFILL_7_DFFSR_18 gnd vdd FILL
XFILL_2_NAND2X1_82 gnd vdd FILL
XFILL_7_DFFSR_29 gnd vdd FILL
XFILL_4_DFFSR_246 gnd vdd FILL
XFILL_33_DFFSR_15 gnd vdd FILL
XFILL_4_DFFSR_257 gnd vdd FILL
XFILL_2_NAND2X1_93 gnd vdd FILL
XFILL_12_BUFX4_100 gnd vdd FILL
XFILL_4_DFFSR_268 gnd vdd FILL
XFILL_33_DFFSR_26 gnd vdd FILL
XFILL_33_DFFSR_37 gnd vdd FILL
XFILL_8_DFFSR_201 gnd vdd FILL
XFILL_33_DFFSR_48 gnd vdd FILL
XFILL_5_NAND3X1_1 gnd vdd FILL
XFILL_10_CLKBUF1_13 gnd vdd FILL
XFILL_8_DFFSR_212 gnd vdd FILL
XFILL_33_DFFSR_59 gnd vdd FILL
XFILL_10_CLKBUF1_24 gnd vdd FILL
XFILL_8_DFFSR_223 gnd vdd FILL
XFILL_8_DFFSR_234 gnd vdd FILL
XFILL_10_CLKBUF1_35 gnd vdd FILL
XFILL_8_DFFSR_245 gnd vdd FILL
XFILL_20_4_2 gnd vdd FILL
XFILL_73_DFFSR_14 gnd vdd FILL
XFILL_8_DFFSR_256 gnd vdd FILL
XFILL_8_DFFSR_267 gnd vdd FILL
XFILL_73_DFFSR_25 gnd vdd FILL
XFILL_73_DFFSR_36 gnd vdd FILL
XFILL_16_MUX2X1_4 gnd vdd FILL
XFILL_73_DFFSR_47 gnd vdd FILL
XFILL_73_DFFSR_58 gnd vdd FILL
XFILL_73_DFFSR_69 gnd vdd FILL
XFILL_42_DFFSR_13 gnd vdd FILL
XFILL_20_DFFSR_200 gnd vdd FILL
XFILL_7_BUFX4_70 gnd vdd FILL
XFILL_42_DFFSR_24 gnd vdd FILL
XFILL_20_DFFSR_211 gnd vdd FILL
XFILL_42_DFFSR_35 gnd vdd FILL
XFILL_7_BUFX4_81 gnd vdd FILL
XFILL_19_MUX2X1_104 gnd vdd FILL
XFILL_10_NOR2X1_13 gnd vdd FILL
XFILL_20_DFFSR_222 gnd vdd FILL
XFILL_7_BUFX4_92 gnd vdd FILL
XFILL_19_MUX2X1_115 gnd vdd FILL
XFILL_42_DFFSR_46 gnd vdd FILL
XFILL_10_NOR2X1_24 gnd vdd FILL
XFILL_1_AOI22X1_7 gnd vdd FILL
XFILL_42_DFFSR_57 gnd vdd FILL
XFILL_20_DFFSR_233 gnd vdd FILL
XFILL_19_MUX2X1_126 gnd vdd FILL
XFILL_10_NOR2X1_35 gnd vdd FILL
XFILL_42_DFFSR_68 gnd vdd FILL
XFILL_19_MUX2X1_137 gnd vdd FILL
XFILL_20_DFFSR_244 gnd vdd FILL
XFILL_10_NOR2X1_46 gnd vdd FILL
XFILL_20_DFFSR_255 gnd vdd FILL
XFILL_19_MUX2X1_148 gnd vdd FILL
XFILL_42_DFFSR_79 gnd vdd FILL
XFILL_10_NOR2X1_57 gnd vdd FILL
XFILL_19_MUX2X1_159 gnd vdd FILL
XFILL_6_AOI21X1_60 gnd vdd FILL
XFILL_20_DFFSR_266 gnd vdd FILL
XFILL_6_AOI21X1_71 gnd vdd FILL
XFILL_10_NOR2X1_68 gnd vdd FILL
XFILL_10_NOR2X1_79 gnd vdd FILL
XFILL_1_INVX1_206 gnd vdd FILL
XFILL_82_DFFSR_12 gnd vdd FILL
XFILL_1_INVX1_217 gnd vdd FILL
XFILL_16_OAI22X1_40 gnd vdd FILL
XFILL_82_DFFSR_23 gnd vdd FILL
XFILL_16_OAI22X1_51 gnd vdd FILL
XFILL_24_DFFSR_210 gnd vdd FILL
XFILL_82_DFFSR_34 gnd vdd FILL
XFILL_24_DFFSR_221 gnd vdd FILL
XFILL_82_DFFSR_45 gnd vdd FILL
XFILL_1_INVX1_228 gnd vdd FILL
XFILL_5_AOI22X1_6 gnd vdd FILL
XFILL_24_DFFSR_232 gnd vdd FILL
XFILL_82_DFFSR_56 gnd vdd FILL
XFILL_11_DFFSR_12 gnd vdd FILL
XFILL_24_DFFSR_243 gnd vdd FILL
XFILL_82_DFFSR_67 gnd vdd FILL
XFILL_11_DFFSR_23 gnd vdd FILL
XFILL_82_DFFSR_78 gnd vdd FILL
XFILL_24_DFFSR_254 gnd vdd FILL
XFILL_11_DFFSR_34 gnd vdd FILL
XFILL_82_DFFSR_89 gnd vdd FILL
XFILL_11_DFFSR_45 gnd vdd FILL
XFILL_24_DFFSR_265 gnd vdd FILL
XFILL_0_CLKBUF1_30 gnd vdd FILL
XFILL_9_NOR2X1_170 gnd vdd FILL
XFILL_0_CLKBUF1_41 gnd vdd FILL
XFILL_11_DFFSR_56 gnd vdd FILL
XFILL_5_INVX1_205 gnd vdd FILL
XFILL_3_5_2 gnd vdd FILL
XFILL_9_NOR2X1_181 gnd vdd FILL
XFILL_28_5_2 gnd vdd FILL
XFILL_11_DFFSR_67 gnd vdd FILL
XFILL_5_INVX1_216 gnd vdd FILL
XFILL_9_NOR2X1_5 gnd vdd FILL
XFILL_51_DFFSR_110 gnd vdd FILL
XFILL_11_DFFSR_78 gnd vdd FILL
XFILL_5_INVX1_227 gnd vdd FILL
XFILL_9_NOR2X1_192 gnd vdd FILL
XFILL_27_0_1 gnd vdd FILL
XFILL_11_DFFSR_89 gnd vdd FILL
XFILL_2_0_1 gnd vdd FILL
XFILL_28_DFFSR_220 gnd vdd FILL
XFILL_51_DFFSR_121 gnd vdd FILL
XFILL_51_DFFSR_132 gnd vdd FILL
XFILL_9_AOI22X1_5 gnd vdd FILL
XFILL_28_DFFSR_231 gnd vdd FILL
XFILL_51_DFFSR_143 gnd vdd FILL
XFILL_28_DFFSR_242 gnd vdd FILL
XFILL_51_DFFSR_11 gnd vdd FILL
XFILL_51_DFFSR_154 gnd vdd FILL
XFILL_51_DFFSR_22 gnd vdd FILL
XFILL_28_DFFSR_253 gnd vdd FILL
XFILL_51_DFFSR_33 gnd vdd FILL
XFILL_2_BUFX2_6 gnd vdd FILL
XFILL_22_NOR3X1_8 gnd vdd FILL
XFILL_51_DFFSR_165 gnd vdd FILL
XFILL_28_DFFSR_264 gnd vdd FILL
XFILL_51_DFFSR_44 gnd vdd FILL
XFILL_28_DFFSR_275 gnd vdd FILL
XFILL_51_DFFSR_55 gnd vdd FILL
XFILL_51_DFFSR_176 gnd vdd FILL
XFILL_51_DFFSR_187 gnd vdd FILL
XFILL_51_DFFSR_198 gnd vdd FILL
XFILL_51_DFFSR_66 gnd vdd FILL
XFILL_51_DFFSR_77 gnd vdd FILL
XFILL_55_DFFSR_120 gnd vdd FILL
XFILL_51_DFFSR_88 gnd vdd FILL
XFILL_55_DFFSR_131 gnd vdd FILL
XFILL_51_DFFSR_99 gnd vdd FILL
XFILL_55_DFFSR_142 gnd vdd FILL
XFILL_55_DFFSR_153 gnd vdd FILL
XFILL_8_MUX2X1_3 gnd vdd FILL
XFILL_55_DFFSR_164 gnd vdd FILL
XFILL_55_DFFSR_175 gnd vdd FILL
XFILL_20_DFFSR_10 gnd vdd FILL
XFILL_55_DFFSR_186 gnd vdd FILL
XFILL_11_4_2 gnd vdd FILL
XFILL_61_DFFSR_5 gnd vdd FILL
XFILL_20_DFFSR_21 gnd vdd FILL
XFILL_55_DFFSR_197 gnd vdd FILL
XFILL_9_MUX2X1_110 gnd vdd FILL
XFILL_9_MUX2X1_121 gnd vdd FILL
XFILL_20_DFFSR_32 gnd vdd FILL
XFILL_20_DFFSR_43 gnd vdd FILL
XFILL_9_MUX2X1_132 gnd vdd FILL
XFILL_59_DFFSR_130 gnd vdd FILL
XFILL_9_MUX2X1_143 gnd vdd FILL
XFILL_20_DFFSR_54 gnd vdd FILL
XFILL_20_DFFSR_65 gnd vdd FILL
XFILL_59_DFFSR_141 gnd vdd FILL
XFILL_59_DFFSR_152 gnd vdd FILL
XFILL_9_MUX2X1_154 gnd vdd FILL
XFILL_20_DFFSR_76 gnd vdd FILL
XFILL_9_MUX2X1_165 gnd vdd FILL
XFILL_59_DFFSR_163 gnd vdd FILL
XFILL_59_DFFSR_174 gnd vdd FILL
XFILL_20_DFFSR_87 gnd vdd FILL
XFILL_9_MUX2X1_176 gnd vdd FILL
XFILL_20_DFFSR_98 gnd vdd FILL
XFILL_2_DFFSR_101 gnd vdd FILL
XFILL_9_MUX2X1_187 gnd vdd FILL
XFILL_5_NOR3X1_9 gnd vdd FILL
XFILL_60_DFFSR_20 gnd vdd FILL
XFILL_2_DFFSR_112 gnd vdd FILL
XFILL_59_DFFSR_185 gnd vdd FILL
XFILL_59_DFFSR_196 gnd vdd FILL
XFILL_60_DFFSR_31 gnd vdd FILL
XFILL_2_DFFSR_123 gnd vdd FILL
XFILL_2_DFFSR_134 gnd vdd FILL
XFILL_31_NOR3X1_6 gnd vdd FILL
XFILL_60_DFFSR_42 gnd vdd FILL
XFILL_2_DFFSR_145 gnd vdd FILL
XFILL_60_DFFSR_53 gnd vdd FILL
XFILL_2_DFFSR_156 gnd vdd FILL
XFILL_60_DFFSR_64 gnd vdd FILL
XFILL_60_DFFSR_75 gnd vdd FILL
XFILL_2_DFFSR_167 gnd vdd FILL
XFILL_2_DFFSR_178 gnd vdd FILL
XFILL_60_DFFSR_86 gnd vdd FILL
XFILL_6_DFFSR_100 gnd vdd FILL
XFILL_2_DFFSR_189 gnd vdd FILL
XFILL_60_DFFSR_97 gnd vdd FILL
XFILL_6_DFFSR_111 gnd vdd FILL
XFILL_37_DFFSR_109 gnd vdd FILL
XFILL_3_DFFSR_11 gnd vdd FILL
XFILL_6_DFFSR_122 gnd vdd FILL
XFILL_10_MUX2X1_20 gnd vdd FILL
XFILL_6_DFFSR_133 gnd vdd FILL
XFILL_3_DFFSR_22 gnd vdd FILL
XFILL_10_MUX2X1_31 gnd vdd FILL
XFILL_6_DFFSR_144 gnd vdd FILL
XFILL_10_MUX2X1_42 gnd vdd FILL
XFILL_3_DFFSR_33 gnd vdd FILL
XFILL_10_MUX2X1_53 gnd vdd FILL
XFILL_6_DFFSR_155 gnd vdd FILL
XFILL_3_DFFSR_44 gnd vdd FILL
XFILL_3_DFFSR_55 gnd vdd FILL
XFILL_10_MUX2X1_64 gnd vdd FILL
XFILL_11_NAND3X1_18 gnd vdd FILL
XFILL_26_DFFSR_8 gnd vdd FILL
XFILL_6_DFFSR_166 gnd vdd FILL
XFILL_3_DFFSR_66 gnd vdd FILL
XFILL_11_NAND3X1_29 gnd vdd FILL
XFILL_83_DFFSR_9 gnd vdd FILL
XFILL_6_DFFSR_177 gnd vdd FILL
XFILL_10_MUX2X1_75 gnd vdd FILL
XFILL_3_DFFSR_77 gnd vdd FILL
XFILL_10_MUX2X1_86 gnd vdd FILL
XFILL_6_DFFSR_188 gnd vdd FILL
XFILL_10_MUX2X1_97 gnd vdd FILL
XFILL_3_DFFSR_88 gnd vdd FILL
XFILL_6_DFFSR_199 gnd vdd FILL
XFILL_3_DFFSR_99 gnd vdd FILL
XFILL_31_CLKBUF1_18 gnd vdd FILL
XFILL_14_MUX2X1_30 gnd vdd FILL
XFILL_31_CLKBUF1_29 gnd vdd FILL
XFILL_14_MUX2X1_41 gnd vdd FILL
XFILL_14_MUX2X1_52 gnd vdd FILL
XFILL_14_MUX2X1_63 gnd vdd FILL
XFILL_19_5_2 gnd vdd FILL
XFILL_14_MUX2X1_74 gnd vdd FILL
XFILL_2_NOR3X1_12 gnd vdd FILL
XFILL_14_MUX2X1_85 gnd vdd FILL
XFILL_2_NOR3X1_23 gnd vdd FILL
XFILL_18_0_1 gnd vdd FILL
XFILL_2_NOR3X1_34 gnd vdd FILL
XFILL_14_MUX2X1_96 gnd vdd FILL
XFILL_2_NOR3X1_45 gnd vdd FILL
XFILL_18_MUX2X1_40 gnd vdd FILL
XFILL_18_MUX2X1_51 gnd vdd FILL
XFILL_61_3_2 gnd vdd FILL
XFILL_0_INVX1_4 gnd vdd FILL
XFILL_18_MUX2X1_62 gnd vdd FILL
XFILL_18_MUX2X1_73 gnd vdd FILL
XFILL_6_NOR3X1_11 gnd vdd FILL
XFILL_18_MUX2X1_84 gnd vdd FILL
XFILL_6_NOR3X1_22 gnd vdd FILL
XFILL_6_NOR3X1_33 gnd vdd FILL
XFILL_18_MUX2X1_95 gnd vdd FILL
XFILL_22_6 gnd vdd FILL
XFILL_6_NOR3X1_44 gnd vdd FILL
XFILL_22_DFFSR_120 gnd vdd FILL
XFILL_15_5 gnd vdd FILL
XFILL_87_DFFSR_209 gnd vdd FILL
XFILL_22_DFFSR_131 gnd vdd FILL
XFILL_30_7_0 gnd vdd FILL
XFILL_22_DFFSR_142 gnd vdd FILL
XFILL_22_DFFSR_153 gnd vdd FILL
XFILL_22_DFFSR_164 gnd vdd FILL
XFILL_3_INVX1_104 gnd vdd FILL
XFILL_22_DFFSR_175 gnd vdd FILL
XFILL_3_INVX1_115 gnd vdd FILL
XFILL_22_DFFSR_186 gnd vdd FILL
XFILL_22_DFFSR_197 gnd vdd FILL
XFILL_3_INVX1_126 gnd vdd FILL
XFILL_3_INVX1_137 gnd vdd FILL
XFILL_1_NAND3X1_13 gnd vdd FILL
XFILL_26_DFFSR_130 gnd vdd FILL
XFILL_3_INVX1_148 gnd vdd FILL
XFILL_1_NAND3X1_24 gnd vdd FILL
XFILL_3_INVX1_159 gnd vdd FILL
XFILL_1_NAND3X1_35 gnd vdd FILL
XFILL_26_DFFSR_141 gnd vdd FILL
XFILL_26_DFFSR_152 gnd vdd FILL
XFILL_1_NAND3X1_46 gnd vdd FILL
XFILL_1_NAND3X1_57 gnd vdd FILL
XFILL_26_DFFSR_163 gnd vdd FILL
XFILL_26_DFFSR_174 gnd vdd FILL
XFILL_5_NAND2X1_15 gnd vdd FILL
XFILL_5_NAND2X1_26 gnd vdd FILL
XFILL_1_NAND3X1_68 gnd vdd FILL
XFILL_7_INVX1_103 gnd vdd FILL
XFILL_7_INVX1_114 gnd vdd FILL
XFILL_1_NAND3X1_79 gnd vdd FILL
XFILL_5_NAND2X1_37 gnd vdd FILL
XFILL_26_DFFSR_185 gnd vdd FILL
XFILL_26_DFFSR_196 gnd vdd FILL
XFILL_7_INVX1_125 gnd vdd FILL
XFILL_5_NAND2X1_48 gnd vdd FILL
XINVX1_150 INVX1_150/A gnd NOR2X1_47/A vdd INVX1
XFILL_5_NAND2X1_59 gnd vdd FILL
XFILL_7_INVX1_136 gnd vdd FILL
XINVX1_161 INVX1_161/A gnd INVX1_161/Y vdd INVX1
XFILL_7_INVX1_147 gnd vdd FILL
XINVX1_172 INVX1_172/A gnd INVX1_172/Y vdd INVX1
XFILL_7_INVX1_158 gnd vdd FILL
XFILL_7_INVX1_169 gnd vdd FILL
XINVX1_183 INVX1_183/A gnd INVX1_183/Y vdd INVX1
XINVX1_194 DFFSR_96/Q gnd INVX1_194/Y vdd INVX1
XFILL_22_NOR3X1_20 gnd vdd FILL
XFILL_22_NOR3X1_31 gnd vdd FILL
XFILL_22_NOR3X1_42 gnd vdd FILL
XFILL_15_MUX2X1_190 gnd vdd FILL
XFILL_72_DFFSR_220 gnd vdd FILL
XFILL_72_DFFSR_231 gnd vdd FILL
XFILL_72_DFFSR_242 gnd vdd FILL
XFILL_72_DFFSR_253 gnd vdd FILL
XFILL_72_DFFSR_264 gnd vdd FILL
XFILL_72_DFFSR_275 gnd vdd FILL
XFILL_26_NOR3X1_30 gnd vdd FILL
XFILL_26_NOR3X1_41 gnd vdd FILL
XFILL_26_NOR3X1_52 gnd vdd FILL
XFILL_76_DFFSR_230 gnd vdd FILL
XFILL_11_NOR2X1_108 gnd vdd FILL
XFILL_5_OAI22X1_9 gnd vdd FILL
XFILL_76_DFFSR_241 gnd vdd FILL
XFILL_11_NOR2X1_119 gnd vdd FILL
XFILL_1_NOR3X1_2 gnd vdd FILL
XFILL_76_DFFSR_252 gnd vdd FILL
XFILL_76_DFFSR_263 gnd vdd FILL
XFILL_76_DFFSR_274 gnd vdd FILL
XFILL_31_CLKBUF1_4 gnd vdd FILL
XFILL_52_3_2 gnd vdd FILL
XFILL_9_AOI21X1_15 gnd vdd FILL
XFILL_9_OAI22X1_8 gnd vdd FILL
XFILL_9_AOI21X1_26 gnd vdd FILL
XFILL_9_AOI21X1_37 gnd vdd FILL
XFILL_9_AOI21X1_48 gnd vdd FILL
XFILL_9_AOI21X1_59 gnd vdd FILL
XFILL_19_OAI22X1_17 gnd vdd FILL
XFILL_21_7_0 gnd vdd FILL
XFILL_35_CLKBUF1_3 gnd vdd FILL
XFILL_19_OAI22X1_28 gnd vdd FILL
XFILL_20_CLKBUF1_14 gnd vdd FILL
XFILL_20_CLKBUF1_25 gnd vdd FILL
XFILL_19_OAI22X1_39 gnd vdd FILL
XFILL_54_DFFSR_209 gnd vdd FILL
XFILL_20_CLKBUF1_36 gnd vdd FILL
XFILL_43_DFFSR_2 gnd vdd FILL
XFILL_3_CLKBUF1_18 gnd vdd FILL
XFILL_3_CLKBUF1_29 gnd vdd FILL
XFILL_81_DFFSR_109 gnd vdd FILL
XFILL_58_DFFSR_208 gnd vdd FILL
XFILL_58_DFFSR_219 gnd vdd FILL
XFILL_6_BUFX2_7 gnd vdd FILL
XFILL_85_DFFSR_108 gnd vdd FILL
XFILL_1_NOR2X1_103 gnd vdd FILL
XFILL_1_NOR2X1_114 gnd vdd FILL
XFILL_85_DFFSR_119 gnd vdd FILL
XFILL_12_OAI21X1_19 gnd vdd FILL
XFILL_1_NOR2X1_125 gnd vdd FILL
XFILL_1_NOR2X1_136 gnd vdd FILL
XFILL_1_NOR2X1_147 gnd vdd FILL
XFILL_1_NOR2X1_158 gnd vdd FILL
XFILL_1_NOR2X1_169 gnd vdd FILL
XFILL_65_DFFSR_6 gnd vdd FILL
XFILL_8_BUFX4_15 gnd vdd FILL
XFILL_8_BUFX4_26 gnd vdd FILL
XFILL_8_BUFX4_37 gnd vdd FILL
XFILL_11_NAND2X1_40 gnd vdd FILL
XFILL_11_NAND2X1_51 gnd vdd FILL
XFILL_11_NAND2X1_62 gnd vdd FILL
XFILL_8_BUFX4_48 gnd vdd FILL
XFILL_11_NAND2X1_73 gnd vdd FILL
XFILL_8_BUFX4_59 gnd vdd FILL
XFILL_9_OAI22X1_12 gnd vdd FILL
XFILL_9_OAI22X1_23 gnd vdd FILL
XFILL_9_OAI22X1_34 gnd vdd FILL
XFILL_11_NAND2X1_84 gnd vdd FILL
XFILL_11_NAND2X1_95 gnd vdd FILL
XFILL_9_OAI22X1_45 gnd vdd FILL
XFILL_43_DFFSR_230 gnd vdd FILL
XFILL_43_3_2 gnd vdd FILL
XFILL_43_DFFSR_241 gnd vdd FILL
XFILL_43_DFFSR_252 gnd vdd FILL
XNAND3X1_103 INVX1_103/A BUFX4_60/Y AND2X2_1/Y gnd NAND3X1_106/A vdd NAND3X1
XFILL_43_DFFSR_263 gnd vdd FILL
XFILL_43_DFFSR_274 gnd vdd FILL
XFILL_1_MUX2X1_109 gnd vdd FILL
XNAND3X1_114 DFFSR_150/Q BUFX4_91/Y NOR3X1_9/Y gnd NAND2X1_69/B vdd NAND3X1
XNAND3X1_125 NAND3X1_125/A NAND3X1_125/B NAND3X1_125/C gnd INVX1_128/A vdd NAND3X1
XFILL_5_BUFX4_1 gnd vdd FILL
XFILL_6_NOR2X1_203 gnd vdd FILL
XFILL_70_DFFSR_130 gnd vdd FILL
XFILL_12_7_0 gnd vdd FILL
XFILL_47_DFFSR_240 gnd vdd FILL
XFILL_70_DFFSR_141 gnd vdd FILL
XFILL_70_DFFSR_152 gnd vdd FILL
XFILL_47_DFFSR_251 gnd vdd FILL
XFILL_70_DFFSR_163 gnd vdd FILL
XFILL_47_DFFSR_262 gnd vdd FILL
XFILL_15_AND2X2_3 gnd vdd FILL
XFILL_70_DFFSR_174 gnd vdd FILL
XFILL_2_OAI21X1_14 gnd vdd FILL
XFILL_47_DFFSR_273 gnd vdd FILL
XFILL_70_DFFSR_185 gnd vdd FILL
XFILL_2_OAI21X1_25 gnd vdd FILL
XFILL_70_DFFSR_196 gnd vdd FILL
XFILL_2_OAI21X1_36 gnd vdd FILL
XFILL_21_DFFSR_209 gnd vdd FILL
XFILL_2_OAI21X1_47 gnd vdd FILL
XFILL_74_DFFSR_140 gnd vdd FILL
XFILL_74_DFFSR_151 gnd vdd FILL
XFILL_74_DFFSR_162 gnd vdd FILL
XFILL_74_DFFSR_173 gnd vdd FILL
XFILL_15_AOI21X1_40 gnd vdd FILL
XFILL_74_DFFSR_184 gnd vdd FILL
XFILL_15_AOI21X1_51 gnd vdd FILL
XFILL_74_DFFSR_195 gnd vdd FILL
XFILL_15_AOI21X1_62 gnd vdd FILL
XFILL_25_DFFSR_208 gnd vdd FILL
XFILL_15_AOI21X1_73 gnd vdd FILL
XFILL_12_BUFX4_20 gnd vdd FILL
XFILL_25_DFFSR_219 gnd vdd FILL
XFILL_4_INVX1_5 gnd vdd FILL
XFILL_12_BUFX4_31 gnd vdd FILL
XFILL_1_NAND2X1_90 gnd vdd FILL
XFILL_12_BUFX4_42 gnd vdd FILL
XFILL_78_DFFSR_150 gnd vdd FILL
XFILL_78_DFFSR_161 gnd vdd FILL
XFILL_12_BUFX4_53 gnd vdd FILL
XFILL_12_BUFX4_64 gnd vdd FILL
XFILL_78_DFFSR_172 gnd vdd FILL
XFILL_78_DFFSR_183 gnd vdd FILL
XFILL_12_BUFX4_75 gnd vdd FILL
XFILL_12_BUFX4_86 gnd vdd FILL
XFILL_52_DFFSR_108 gnd vdd FILL
XFILL_78_DFFSR_194 gnd vdd FILL
XFILL_29_DFFSR_207 gnd vdd FILL
XFILL_12_BUFX4_97 gnd vdd FILL
XFILL_52_DFFSR_119 gnd vdd FILL
XFILL_29_DFFSR_218 gnd vdd FILL
XFILL_29_DFFSR_229 gnd vdd FILL
XFILL_56_DFFSR_107 gnd vdd FILL
XFILL_56_DFFSR_118 gnd vdd FILL
XFILL_56_DFFSR_129 gnd vdd FILL
XFILL_5_INVX4_1 gnd vdd FILL
XFILL_62_6_0 gnd vdd FILL
XFILL_30_DFFSR_19 gnd vdd FILL
XFILL_6_INVX1_10 gnd vdd FILL
XFILL_34_3_2 gnd vdd FILL
XFILL_6_INVX1_21 gnd vdd FILL
XFILL_6_INVX1_32 gnd vdd FILL
XFILL_18_MUX2X1_101 gnd vdd FILL
XFILL_18_MUX2X1_112 gnd vdd FILL
XFILL_6_INVX1_43 gnd vdd FILL
XFILL_7_AND2X2_2 gnd vdd FILL
XFILL_18_MUX2X1_123 gnd vdd FILL
XFILL_10_DFFSR_230 gnd vdd FILL
XFILL_6_INVX1_54 gnd vdd FILL
XFILL_6_INVX1_65 gnd vdd FILL
XFILL_20_3 gnd vdd FILL
XFILL_10_DFFSR_241 gnd vdd FILL
XFILL_18_MUX2X1_134 gnd vdd FILL
XFILL_18_MUX2X1_145 gnd vdd FILL
XFILL_10_DFFSR_252 gnd vdd FILL
XFILL_6_INVX1_76 gnd vdd FILL
XFILL_18_MUX2X1_156 gnd vdd FILL
XFILL_6_INVX1_87 gnd vdd FILL
XFILL_10_DFFSR_263 gnd vdd FILL
XFILL_10_DFFSR_274 gnd vdd FILL
XFILL_6_INVX1_98 gnd vdd FILL
XFILL_18_MUX2X1_167 gnd vdd FILL
XFILL_70_DFFSR_18 gnd vdd FILL
XFILL_70_DFFSR_29 gnd vdd FILL
XFILL_18_MUX2X1_178 gnd vdd FILL
XFILL_13_2 gnd vdd FILL
XFILL_18_MUX2X1_189 gnd vdd FILL
XFILL_13_MUX2X1_8 gnd vdd FILL
XFILL_14_DFFSR_240 gnd vdd FILL
XDFFSR_101 INVX1_105/A DFFSR_57/CLK BUFX4_21/Y vdd MUX2X1_92/Y gnd vdd DFFSR
XFILL_14_DFFSR_251 gnd vdd FILL
XFILL_14_DFFSR_262 gnd vdd FILL
XDFFSR_112 INVX2_5/A CLKBUF1_24/Y BUFX4_32/Y vdd DFFSR_112/D gnd vdd DFFSR
XFILL_7_DFFSR_109 gnd vdd FILL
XFILL_14_DFFSR_273 gnd vdd FILL
XDFFSR_123 INVX1_177/A CLKBUF1_34/Y BUFX4_23/Y vdd DFFSR_123/D gnd vdd DFFSR
XDFFSR_134 INVX1_159/A CLKBUF1_1/Y DFFSR_89/R vdd DFFSR_134/D gnd vdd DFFSR
XFILL_4_BUFX4_30 gnd vdd FILL
XFILL_4_BUFX4_41 gnd vdd FILL
XFILL_11_MUX2X1_18 gnd vdd FILL
XDFFSR_145 INVX1_157/A DFFSR_72/CLK DFFSR_96/R vdd DFFSR_145/D gnd vdd DFFSR
XFILL_11_MUX2X1_29 gnd vdd FILL
XFILL_4_BUFX4_52 gnd vdd FILL
XDFFSR_156 NOR2X1_79/A DFFSR_94/CLK DFFSR_98/R vdd DFFSR_156/D gnd vdd DFFSR
XFILL_4_BUFX4_63 gnd vdd FILL
XFILL_2_AOI21X1_5 gnd vdd FILL
XDFFSR_167 NOR2X1_46/A DFFSR_56/CLK DFFSR_56/R vdd DFFSR_167/D gnd vdd DFFSR
XDFFSR_178 INVX1_152/A DFFSR_76/CLK DFFSR_53/R vdd DFFSR_178/D gnd vdd DFFSR
XFILL_41_DFFSR_140 gnd vdd FILL
XFILL_4_BUFX4_74 gnd vdd FILL
XBUFX4_8 BUFX4_8/A gnd BUFX4_8/Y vdd BUFX4
XFILL_4_BUFX4_85 gnd vdd FILL
XFILL_41_DFFSR_151 gnd vdd FILL
XDFFSR_189 INVX1_134/A CLKBUF1_24/Y BUFX4_32/Y vdd INVX1_137/A gnd vdd DFFSR
XFILL_41_DFFSR_162 gnd vdd FILL
XFILL_4_BUFX4_96 gnd vdd FILL
XFILL_18_DFFSR_250 gnd vdd FILL
XFILL_18_DFFSR_261 gnd vdd FILL
XFILL_18_DFFSR_272 gnd vdd FILL
XFILL_41_DFFSR_173 gnd vdd FILL
XFILL_41_DFFSR_184 gnd vdd FILL
XFILL_15_MUX2X1_17 gnd vdd FILL
XFILL_41_DFFSR_195 gnd vdd FILL
XFILL_15_MUX2X1_28 gnd vdd FILL
XFILL_15_MUX2X1_39 gnd vdd FILL
XFILL_6_AOI21X1_4 gnd vdd FILL
XFILL_45_DFFSR_150 gnd vdd FILL
XFILL_45_DFFSR_161 gnd vdd FILL
XFILL_45_DFFSR_172 gnd vdd FILL
XFILL_22_MUX2X1_6 gnd vdd FILL
XFILL_45_DFFSR_183 gnd vdd FILL
XFILL_19_MUX2X1_16 gnd vdd FILL
XFILL_45_DFFSR_194 gnd vdd FILL
XFILL_19_MUX2X1_27 gnd vdd FILL
XFILL_47_DFFSR_3 gnd vdd FILL
XFILL_19_MUX2X1_38 gnd vdd FILL
XFILL_8_MUX2X1_140 gnd vdd FILL
XFILL_19_MUX2X1_49 gnd vdd FILL
XFILL_6_NOR2X1_9 gnd vdd FILL
XNOR3X1_12 INVX1_63/Y NOR3X1_39/C INVX2_2/Y gnd NOR3X1_23/B vdd NOR3X1
XFILL_11_AOI22X1_1 gnd vdd FILL
XFILL_8_MUX2X1_151 gnd vdd FILL
XFILL_49_DFFSR_160 gnd vdd FILL
XFILL_8_MUX2X1_162 gnd vdd FILL
XNOR3X1_23 NOR3X1_1/Y NOR3X1_23/B OAI22X1_1/Y gnd NOR3X1_23/Y vdd NOR3X1
XNOR3X1_34 INVX1_46/Y NOR3X1_49/B NOR3X1_39/C gnd NOR3X1_50/B vdd NOR3X1
XFILL_8_MUX2X1_173 gnd vdd FILL
XFILL_49_DFFSR_171 gnd vdd FILL
XFILL_8_MUX2X1_184 gnd vdd FILL
XFILL_49_DFFSR_182 gnd vdd FILL
XNOR3X1_45 NOR3X1_45/A NOR3X1_49/B NOR3X1_1/B gnd NOR3X1_50/A vdd NOR3X1
XFILL_23_DFFSR_107 gnd vdd FILL
XFILL_49_DFFSR_193 gnd vdd FILL
XFILL_23_DFFSR_118 gnd vdd FILL
XFILL_23_DFFSR_129 gnd vdd FILL
XFILL_53_6_0 gnd vdd FILL
XFILL_0_3_2 gnd vdd FILL
XFILL_25_3_2 gnd vdd FILL
XFILL_5_MUX2X1_7 gnd vdd FILL
XFILL_27_DFFSR_106 gnd vdd FILL
XFILL_27_DFFSR_117 gnd vdd FILL
XFILL_27_DFFSR_128 gnd vdd FILL
XFILL_31_DFFSR_9 gnd vdd FILL
XFILL_27_DFFSR_139 gnd vdd FILL
XFILL_10_NAND3X1_15 gnd vdd FILL
XFILL_10_NAND3X1_26 gnd vdd FILL
XFILL_10_NAND3X1_37 gnd vdd FILL
XFILL_10_NAND3X1_48 gnd vdd FILL
XFILL_69_DFFSR_7 gnd vdd FILL
XFILL_10_NAND3X1_59 gnd vdd FILL
XFILL_30_CLKBUF1_15 gnd vdd FILL
XFILL_39_DFFSR_30 gnd vdd FILL
XFILL_30_CLKBUF1_26 gnd vdd FILL
XFILL_39_DFFSR_41 gnd vdd FILL
XFILL_30_CLKBUF1_37 gnd vdd FILL
XFILL_39_DFFSR_52 gnd vdd FILL
XFILL_39_DFFSR_63 gnd vdd FILL
XFILL_39_DFFSR_74 gnd vdd FILL
XFILL_39_DFFSR_85 gnd vdd FILL
XFILL_23_NOR3X1_18 gnd vdd FILL
XFILL_39_DFFSR_96 gnd vdd FILL
XFILL_23_NOR3X1_29 gnd vdd FILL
XFILL_73_DFFSR_207 gnd vdd FILL
XFILL_79_DFFSR_40 gnd vdd FILL
XFILL_73_DFFSR_218 gnd vdd FILL
XFILL_0_DFFSR_15 gnd vdd FILL
XFILL_79_DFFSR_51 gnd vdd FILL
XFILL_73_DFFSR_229 gnd vdd FILL
XFILL_10_NOR2X1_3 gnd vdd FILL
XFILL_0_DFFSR_26 gnd vdd FILL
XFILL_79_DFFSR_62 gnd vdd FILL
XFILL_0_DFFSR_37 gnd vdd FILL
XFILL_79_DFFSR_73 gnd vdd FILL
XFILL_79_DFFSR_84 gnd vdd FILL
XFILL_0_DFFSR_48 gnd vdd FILL
XFILL_79_DFFSR_95 gnd vdd FILL
XFILL_27_NOR3X1_17 gnd vdd FILL
XFILL_0_DFFSR_59 gnd vdd FILL
XFILL_27_NOR3X1_28 gnd vdd FILL
XFILL_27_NOR3X1_39 gnd vdd FILL
XFILL_9_BUFX4_2 gnd vdd FILL
XFILL_8_4_2 gnd vdd FILL
XFILL_77_DFFSR_206 gnd vdd FILL
XFILL_77_DFFSR_217 gnd vdd FILL
XFILL_2_INVX1_80 gnd vdd FILL
XFILL_77_DFFSR_228 gnd vdd FILL
XFILL_12_DFFSR_150 gnd vdd FILL
XFILL_77_DFFSR_239 gnd vdd FILL
XFILL_12_DFFSR_161 gnd vdd FILL
XFILL_2_INVX1_91 gnd vdd FILL
XFILL_19_NOR3X1_3 gnd vdd FILL
XFILL_12_DFFSR_172 gnd vdd FILL
XFILL_1_CLKBUF1_4 gnd vdd FILL
XFILL_48_DFFSR_50 gnd vdd FILL
XFILL_12_DFFSR_183 gnd vdd FILL
XFILL_12_DFFSR_194 gnd vdd FILL
XFILL_48_DFFSR_61 gnd vdd FILL
XFILL_0_NAND3X1_10 gnd vdd FILL
XFILL_48_DFFSR_72 gnd vdd FILL
XFILL_48_DFFSR_83 gnd vdd FILL
XFILL_0_NAND3X1_21 gnd vdd FILL
XFILL_48_DFFSR_94 gnd vdd FILL
XFILL_0_NAND3X1_32 gnd vdd FILL
XFILL_0_NAND3X1_43 gnd vdd FILL
XFILL_16_DFFSR_160 gnd vdd FILL
XFILL_0_NAND3X1_54 gnd vdd FILL
XFILL_0_NAND3X1_65 gnd vdd FILL
XFILL_5_CLKBUF1_3 gnd vdd FILL
XFILL_4_NAND2X1_12 gnd vdd FILL
XFILL_16_DFFSR_171 gnd vdd FILL
XFILL_4_NAND2X1_23 gnd vdd FILL
XFILL_16_DFFSR_182 gnd vdd FILL
XFILL_0_NAND3X1_76 gnd vdd FILL
XFILL_4_NAND2X1_34 gnd vdd FILL
XFILL_44_6_0 gnd vdd FILL
XFILL_0_NAND3X1_87 gnd vdd FILL
XFILL_16_DFFSR_193 gnd vdd FILL
XFILL_4_NAND2X1_45 gnd vdd FILL
XFILL_16_3_2 gnd vdd FILL
XFILL_0_NAND3X1_98 gnd vdd FILL
XFILL_4_NAND2X1_56 gnd vdd FILL
XFILL_4_NAND2X1_67 gnd vdd FILL
XFILL_4_NAND2X1_78 gnd vdd FILL
XFILL_17_DFFSR_60 gnd vdd FILL
XFILL_4_NAND2X1_89 gnd vdd FILL
XFILL_17_DFFSR_71 gnd vdd FILL
XFILL_17_DFFSR_82 gnd vdd FILL
XFILL_9_CLKBUF1_2 gnd vdd FILL
XFILL_17_DFFSR_93 gnd vdd FILL
XFILL_28_NOR3X1_1 gnd vdd FILL
XFILL_12_NOR3X1_50 gnd vdd FILL
XFILL_57_DFFSR_70 gnd vdd FILL
XFILL_57_DFFSR_81 gnd vdd FILL
XFILL_57_DFFSR_92 gnd vdd FILL
XFILL_62_DFFSR_250 gnd vdd FILL
XFILL_62_DFFSR_261 gnd vdd FILL
XFILL_62_DFFSR_272 gnd vdd FILL
XFILL_2_NOR2X1_2 gnd vdd FILL
XFILL_10_NOR2X1_105 gnd vdd FILL
XFILL_10_NOR2X1_116 gnd vdd FILL
XFILL_10_NOR2X1_127 gnd vdd FILL
XFILL_4_AOI22X1_10 gnd vdd FILL
XFILL_10_NOR2X1_138 gnd vdd FILL
XFILL_10_NOR2X1_149 gnd vdd FILL
XFILL_66_DFFSR_260 gnd vdd FILL
XFILL_66_DFFSR_271 gnd vdd FILL
XFILL_21_CLKBUF1_1 gnd vdd FILL
XFILL_26_DFFSR_80 gnd vdd FILL
XFILL_40_DFFSR_207 gnd vdd FILL
XFILL_26_DFFSR_91 gnd vdd FILL
XFILL_8_AOI21X1_12 gnd vdd FILL
XFILL_40_DFFSR_218 gnd vdd FILL
XFILL_2_OAI21X1_8 gnd vdd FILL
XFILL_40_DFFSR_229 gnd vdd FILL
XFILL_8_AOI21X1_23 gnd vdd FILL
XFILL_8_AOI21X1_34 gnd vdd FILL
XFILL_8_AOI21X1_45 gnd vdd FILL
XFILL_18_OAI22X1_14 gnd vdd FILL
XFILL_8_AOI21X1_56 gnd vdd FILL
XFILL_8_AOI21X1_67 gnd vdd FILL
XFILL_18_OAI22X1_25 gnd vdd FILL
XFILL_8_AOI21X1_78 gnd vdd FILL
XFILL_66_DFFSR_90 gnd vdd FILL
XFILL_18_OAI22X1_36 gnd vdd FILL
XFILL_3_NOR2X1_10 gnd vdd FILL
XFILL_44_DFFSR_206 gnd vdd FILL
XFILL_18_OAI22X1_47 gnd vdd FILL
XFILL_3_NOR2X1_21 gnd vdd FILL
XFILL_44_DFFSR_217 gnd vdd FILL
XFILL_3_NOR2X1_32 gnd vdd FILL
XFILL_6_OAI21X1_7 gnd vdd FILL
XFILL_44_DFFSR_228 gnd vdd FILL
XFILL_3_NOR2X1_43 gnd vdd FILL
XFILL_44_DFFSR_239 gnd vdd FILL
XFILL_66_2_2 gnd vdd FILL
XFILL_3_NOR2X1_54 gnd vdd FILL
XFILL_3_NOR2X1_65 gnd vdd FILL
XFILL_3_NOR2X1_76 gnd vdd FILL
XFILL_86_DFFSR_1 gnd vdd FILL
XFILL_2_CLKBUF1_15 gnd vdd FILL
XFILL_2_CLKBUF1_26 gnd vdd FILL
XFILL_3_NOR2X1_87 gnd vdd FILL
XFILL_2_CLKBUF1_37 gnd vdd FILL
XFILL_71_DFFSR_106 gnd vdd FILL
XFILL_3_NOR2X1_98 gnd vdd FILL
XFILL_9_DFFSR_70 gnd vdd FILL
XFILL_48_DFFSR_205 gnd vdd FILL
XFILL_71_DFFSR_117 gnd vdd FILL
XFILL_7_NOR2X1_20 gnd vdd FILL
XFILL_9_DFFSR_81 gnd vdd FILL
XFILL_7_NOR2X1_31 gnd vdd FILL
XFILL_48_DFFSR_216 gnd vdd FILL
XFILL_9_DFFSR_92 gnd vdd FILL
XFILL_48_DFFSR_227 gnd vdd FILL
XFILL_71_DFFSR_128 gnd vdd FILL
XFILL_7_NOR2X1_42 gnd vdd FILL
XFILL_35_6_0 gnd vdd FILL
XFILL_48_DFFSR_238 gnd vdd FILL
XFILL_71_DFFSR_139 gnd vdd FILL
XFILL_7_NOR2X1_53 gnd vdd FILL
XFILL_11_OAI22X1_4 gnd vdd FILL
XFILL_48_DFFSR_249 gnd vdd FILL
XFILL_7_NOR2X1_64 gnd vdd FILL
XFILL_7_NOR2X1_75 gnd vdd FILL
XFILL_7_NOR2X1_86 gnd vdd FILL
XFILL_75_DFFSR_105 gnd vdd FILL
XFILL_7_NOR2X1_97 gnd vdd FILL
XFILL_0_NOR2X1_100 gnd vdd FILL
XFILL_0_NOR2X1_111 gnd vdd FILL
XFILL_75_DFFSR_116 gnd vdd FILL
XFILL_11_OAI21X1_16 gnd vdd FILL
XFILL_75_DFFSR_127 gnd vdd FILL
XFILL_0_NOR2X1_122 gnd vdd FILL
XFILL_11_OAI21X1_27 gnd vdd FILL
XFILL_75_DFFSR_138 gnd vdd FILL
XFILL_0_DFFSR_8 gnd vdd FILL
XFILL_0_NOR2X1_133 gnd vdd FILL
XFILL_11_OAI21X1_38 gnd vdd FILL
XFILL_75_DFFSR_149 gnd vdd FILL
XFILL_11_OAI21X1_49 gnd vdd FILL
XFILL_15_OAI22X1_3 gnd vdd FILL
XFILL_0_NOR2X1_144 gnd vdd FILL
XFILL_13_DFFSR_6 gnd vdd FILL
XFILL_0_NOR2X1_155 gnd vdd FILL
XFILL_0_NOR2X1_166 gnd vdd FILL
XFILL_0_NOR2X1_177 gnd vdd FILL
XFILL_70_DFFSR_7 gnd vdd FILL
XFILL_79_DFFSR_104 gnd vdd FILL
XFILL_0_NOR2X1_188 gnd vdd FILL
XFILL_0_NOR2X1_199 gnd vdd FILL
XFILL_79_DFFSR_115 gnd vdd FILL
XFILL_79_DFFSR_126 gnd vdd FILL
XFILL_79_DFFSR_137 gnd vdd FILL
XFILL_19_OAI22X1_2 gnd vdd FILL
XFILL_79_DFFSR_148 gnd vdd FILL
XFILL_10_NAND2X1_70 gnd vdd FILL
XFILL_10_NAND2X1_81 gnd vdd FILL
XFILL_8_OAI22X1_20 gnd vdd FILL
XFILL_79_DFFSR_159 gnd vdd FILL
XFILL_8_OAI22X1_31 gnd vdd FILL
XFILL_8_OAI22X1_42 gnd vdd FILL
XFILL_10_NAND2X1_92 gnd vdd FILL
XBUFX2_5 INVX2_5/A gnd addr[1] vdd BUFX2
XFILL_33_DFFSR_260 gnd vdd FILL
XFILL_33_DFFSR_271 gnd vdd FILL
XFILL_0_MUX2X1_106 gnd vdd FILL
XFILL_0_MUX2X1_117 gnd vdd FILL
XFILL_3_NAND2X1_9 gnd vdd FILL
XFILL_0_MUX2X1_128 gnd vdd FILL
XFILL_5_NOR2X1_200 gnd vdd FILL
XFILL_0_MUX2X1_139 gnd vdd FILL
XFILL_5_BUFX4_19 gnd vdd FILL
XFILL_60_DFFSR_160 gnd vdd FILL
XFILL_60_DFFSR_171 gnd vdd FILL
XFILL_1_OAI21X1_11 gnd vdd FILL
XFILL_37_DFFSR_270 gnd vdd FILL
XFILL_1_OAI21X1_22 gnd vdd FILL
XFILL_60_DFFSR_182 gnd vdd FILL
XFILL_7_NAND2X1_8 gnd vdd FILL
XFILL_57_2_2 gnd vdd FILL
XFILL_60_DFFSR_193 gnd vdd FILL
XFILL_11_DFFSR_206 gnd vdd FILL
XFILL_1_OAI21X1_33 gnd vdd FILL
XFILL_11_DFFSR_217 gnd vdd FILL
XFILL_1_OAI21X1_44 gnd vdd FILL
XFILL_3_MUX2X1_50 gnd vdd FILL
XFILL_11_DFFSR_228 gnd vdd FILL
XFILL_3_MUX2X1_61 gnd vdd FILL
XFILL_19_CLKBUF1_40 gnd vdd FILL
XFILL_3_MUX2X1_72 gnd vdd FILL
XFILL_3_MUX2X1_83 gnd vdd FILL
XFILL_11_DFFSR_239 gnd vdd FILL
XFILL_64_DFFSR_170 gnd vdd FILL
XFILL_3_MUX2X1_94 gnd vdd FILL
XFILL_64_DFFSR_181 gnd vdd FILL
XFILL_26_6_0 gnd vdd FILL
XFILL_1_6_0 gnd vdd FILL
XFILL_64_DFFSR_192 gnd vdd FILL
XFILL_14_AOI21X1_70 gnd vdd FILL
XFILL_15_DFFSR_205 gnd vdd FILL
XFILL_12_NAND3X1_5 gnd vdd FILL
XFILL_14_AOI21X1_81 gnd vdd FILL
XFILL_15_DFFSR_216 gnd vdd FILL
XFILL_15_DFFSR_227 gnd vdd FILL
XFILL_7_MUX2X1_60 gnd vdd FILL
XFILL_7_MUX2X1_71 gnd vdd FILL
XFILL_15_DFFSR_238 gnd vdd FILL
XFILL_7_MUX2X1_82 gnd vdd FILL
XFILL_7_MUX2X1_93 gnd vdd FILL
XFILL_15_DFFSR_249 gnd vdd FILL
XFILL_68_DFFSR_180 gnd vdd FILL
XNOR2X1_190 DFFSR_22/Q NOR2X1_190/B gnd NOR2X1_190/Y vdd NOR2X1
XFILL_68_DFFSR_191 gnd vdd FILL
XFILL_42_DFFSR_105 gnd vdd FILL
XFILL_40_1_2 gnd vdd FILL
XFILL_42_DFFSR_116 gnd vdd FILL
XFILL_12_AND2X2_7 gnd vdd FILL
XFILL_19_DFFSR_204 gnd vdd FILL
XFILL_19_DFFSR_215 gnd vdd FILL
XFILL_42_DFFSR_127 gnd vdd FILL
XFILL_19_DFFSR_226 gnd vdd FILL
XFILL_42_DFFSR_138 gnd vdd FILL
XFILL_19_DFFSR_237 gnd vdd FILL
XINVX2_5 INVX2_5/A gnd INVX2_5/Y vdd INVX2
XFILL_42_DFFSR_149 gnd vdd FILL
XFILL_19_DFFSR_248 gnd vdd FILL
XFILL_19_DFFSR_259 gnd vdd FILL
XFILL_46_DFFSR_104 gnd vdd FILL
XAOI21X1_5 BUFX4_68/Y AOI21X1_7/B AOI21X1_5/C gnd DFFSR_140/D vdd AOI21X1
XFILL_46_DFFSR_115 gnd vdd FILL
XFILL_46_DFFSR_126 gnd vdd FILL
XFILL_46_DFFSR_137 gnd vdd FILL
XFILL_46_DFFSR_148 gnd vdd FILL
XFILL_46_DFFSR_159 gnd vdd FILL
XMUX2X1_130 INVX1_173/Y MUX2X1_7/B NAND2X1_89/Y gnd DFFSR_129/D vdd MUX2X1
XMUX2X1_141 INVX1_184/Y BUFX4_66/Y NAND3X1_1/Y gnd DFFSR_114/D vdd MUX2X1
XMUX2X1_152 BUFX4_98/Y INVX1_195/Y NOR2X1_154/Y gnd DFFSR_97/D vdd MUX2X1
XMUX2X1_163 BUFX4_67/Y INVX1_208/Y NOR2X1_162/Y gnd DFFSR_77/D vdd MUX2X1
XFILL_17_MUX2X1_120 gnd vdd FILL
XFILL_17_MUX2X1_131 gnd vdd FILL
XMUX2X1_174 BUFX4_98/Y INVX1_219/Y NOR2X1_165/Y gnd DFFSR_71/D vdd MUX2X1
XMUX2X1_185 BUFX4_68/Y INVX1_4/Y NOR2X1_168/Y gnd DFFSR_55/D vdd MUX2X1
XFILL_9_7_0 gnd vdd FILL
XFILL_23_MUX2X1_80 gnd vdd FILL
XFILL_17_MUX2X1_142 gnd vdd FILL
XFILL_17_MUX2X1_153 gnd vdd FILL
XFILL_23_MUX2X1_91 gnd vdd FILL
XFILL_17_MUX2X1_164 gnd vdd FILL
XFILL_17_MUX2X1_175 gnd vdd FILL
XFILL_17_MUX2X1_186 gnd vdd FILL
XFILL_16_AOI22X1_9 gnd vdd FILL
XFILL_48_2_2 gnd vdd FILL
XINVX1_70 INVX1_70/A gnd INVX1_70/Y vdd INVX1
XINVX1_81 INVX1_81/A gnd INVX1_81/Y vdd INVX1
XFILL_54_9 gnd vdd FILL
XINVX1_92 INVX1_92/A gnd INVX1_92/Y vdd INVX1
XFILL_3_INVX1_14 gnd vdd FILL
XFILL_10_INVX8_4 gnd vdd FILL
XFILL_3_INVX1_25 gnd vdd FILL
XFILL_3_INVX1_36 gnd vdd FILL
XFILL_17_6_0 gnd vdd FILL
XFILL_3_INVX1_47 gnd vdd FILL
XFILL_4_AND2X2_6 gnd vdd FILL
XFILL_31_DFFSR_170 gnd vdd FILL
XFILL_3_INVX1_58 gnd vdd FILL
XFILL_3_INVX1_69 gnd vdd FILL
XFILL_31_DFFSR_181 gnd vdd FILL
XFILL_49_DFFSR_17 gnd vdd FILL
XFILL_31_DFFSR_192 gnd vdd FILL
XFILL_49_DFFSR_28 gnd vdd FILL
XFILL_49_DFFSR_39 gnd vdd FILL
XFILL_31_1_2 gnd vdd FILL
XFILL_35_DFFSR_180 gnd vdd FILL
XFILL_35_DFFSR_191 gnd vdd FILL
XFILL_1_BUFX4_12 gnd vdd FILL
XFILL_52_DFFSR_4 gnd vdd FILL
XFILL_1_BUFX4_23 gnd vdd FILL
XFILL_1_BUFX4_34 gnd vdd FILL
XFILL_1_BUFX4_45 gnd vdd FILL
XFILL_18_DFFSR_16 gnd vdd FILL
XFILL_1_BUFX4_56 gnd vdd FILL
XFILL_18_DFFSR_27 gnd vdd FILL
XFILL_7_MUX2X1_170 gnd vdd FILL
XFILL_18_DFFSR_38 gnd vdd FILL
XFILL_1_BUFX4_67 gnd vdd FILL
XFILL_1_BUFX4_78 gnd vdd FILL
XFILL_18_DFFSR_49 gnd vdd FILL
XFILL_7_MUX2X1_181 gnd vdd FILL
XFILL_39_DFFSR_190 gnd vdd FILL
XFILL_7_MUX2X1_192 gnd vdd FILL
XFILL_1_BUFX4_89 gnd vdd FILL
XFILL_13_DFFSR_104 gnd vdd FILL
XFILL_13_DFFSR_115 gnd vdd FILL
XFILL_13_DFFSR_126 gnd vdd FILL
XFILL_13_DFFSR_137 gnd vdd FILL
XNOR2X1_3 NOR2X1_3/A NOR2X1_6/B gnd NOR2X1_3/Y vdd NOR2X1
XFILL_13_DFFSR_148 gnd vdd FILL
XFILL_58_DFFSR_15 gnd vdd FILL
XFILL_58_DFFSR_26 gnd vdd FILL
XFILL_13_DFFSR_159 gnd vdd FILL
XFILL_58_DFFSR_37 gnd vdd FILL
XFILL_58_DFFSR_48 gnd vdd FILL
XFILL_58_DFFSR_59 gnd vdd FILL
XFILL_81_DFFSR_270 gnd vdd FILL
XFILL_17_DFFSR_103 gnd vdd FILL
XFILL_17_DFFSR_114 gnd vdd FILL
XFILL_17_DFFSR_125 gnd vdd FILL
XFILL_17_DFFSR_136 gnd vdd FILL
XFILL_4_DFFSR_9 gnd vdd FILL
XFILL_17_DFFSR_147 gnd vdd FILL
XFILL_17_DFFSR_158 gnd vdd FILL
XFILL_17_DFFSR_169 gnd vdd FILL
XFILL_17_DFFSR_7 gnd vdd FILL
XFILL_74_DFFSR_8 gnd vdd FILL
XFILL_27_DFFSR_14 gnd vdd FILL
XFILL_27_DFFSR_25 gnd vdd FILL
XFILL_27_DFFSR_36 gnd vdd FILL
XFILL_39_2_2 gnd vdd FILL
XFILL_27_DFFSR_47 gnd vdd FILL
XFILL_27_DFFSR_58 gnd vdd FILL
XFILL_27_DFFSR_69 gnd vdd FILL
XFILL_67_DFFSR_13 gnd vdd FILL
XFILL_13_NOR3X1_15 gnd vdd FILL
XFILL_13_NOR3X1_26 gnd vdd FILL
XFILL_67_DFFSR_24 gnd vdd FILL
XFILL_13_NOR3X1_37 gnd vdd FILL
XFILL_67_DFFSR_35 gnd vdd FILL
XFILL_13_NOR3X1_48 gnd vdd FILL
XFILL_67_DFFSR_46 gnd vdd FILL
XFILL_63_DFFSR_204 gnd vdd FILL
XFILL_63_DFFSR_215 gnd vdd FILL
XFILL_67_DFFSR_57 gnd vdd FILL
XFILL_67_DFFSR_68 gnd vdd FILL
XFILL_63_DFFSR_226 gnd vdd FILL
XFILL_63_DFFSR_237 gnd vdd FILL
XFILL_67_DFFSR_79 gnd vdd FILL
XFILL_63_DFFSR_248 gnd vdd FILL
XFILL_17_NOR3X1_14 gnd vdd FILL
XFILL_63_DFFSR_259 gnd vdd FILL
XFILL_17_NOR3X1_25 gnd vdd FILL
XFILL_50_4_0 gnd vdd FILL
XFILL_17_NOR3X1_36 gnd vdd FILL
XFILL_17_NOR3X1_47 gnd vdd FILL
XFILL_22_1_2 gnd vdd FILL
XFILL_67_DFFSR_203 gnd vdd FILL
XFILL_36_DFFSR_12 gnd vdd FILL
XFILL_67_DFFSR_214 gnd vdd FILL
XFILL_36_DFFSR_23 gnd vdd FILL
XFILL_67_DFFSR_225 gnd vdd FILL
XFILL_0_OAI22X1_19 gnd vdd FILL
XFILL_67_DFFSR_236 gnd vdd FILL
XFILL_36_DFFSR_34 gnd vdd FILL
XFILL_67_DFFSR_247 gnd vdd FILL
XFILL_36_DFFSR_45 gnd vdd FILL
XFILL_36_DFFSR_56 gnd vdd FILL
XFILL_67_DFFSR_258 gnd vdd FILL
XFILL_67_DFFSR_269 gnd vdd FILL
XFILL_36_DFFSR_67 gnd vdd FILL
XFILL_36_DFFSR_78 gnd vdd FILL
XFILL_36_DFFSR_89 gnd vdd FILL
XAOI21X1_13 BUFX4_81/Y NOR2X1_153/B NOR2X1_149/Y gnd DFFSR_98/D vdd AOI21X1
XAOI21X1_24 BUFX4_83/Y NOR2X1_181/B NOR2X1_178/Y gnd DFFSR_28/D vdd AOI21X1
XFILL_76_DFFSR_11 gnd vdd FILL
XAOI21X1_35 BUFX4_83/Y NOR2X1_195/B NOR2X1_192/Y gnd DFFSR_15/D vdd AOI21X1
XFILL_76_DFFSR_22 gnd vdd FILL
XAOI21X1_46 BUFX4_85/Y NOR2X1_6/B NOR2X1_3/Y gnd DFFSR_271/D vdd AOI21X1
XFILL_76_DFFSR_33 gnd vdd FILL
XAOI21X1_57 MUX2X1_8/A NOR2X1_19/B NOR2X1_18/Y gnd DFFSR_253/D vdd AOI21X1
XFILL_76_DFFSR_44 gnd vdd FILL
XFILL_19_MUX2X1_1 gnd vdd FILL
XAOI21X1_68 DFFSR_6/Q NOR2X1_52/Y NOR2X1_51/Y gnd NAND3X1_55/B vdd AOI21X1
XFILL_76_DFFSR_55 gnd vdd FILL
XAOI21X1_79 OAI21X1_39/Y OAI21X1_40/Y INVX2_3/A gnd OAI21X1_47/A vdd AOI21X1
XFILL_3_NAND2X1_20 gnd vdd FILL
XFILL_76_DFFSR_66 gnd vdd FILL
XFILL_3_NAND2X1_31 gnd vdd FILL
XFILL_76_DFFSR_77 gnd vdd FILL
XFILL_26_CLKBUF1_9 gnd vdd FILL
XFILL_3_NAND2X1_42 gnd vdd FILL
XFILL_76_DFFSR_88 gnd vdd FILL
XFILL_4_NOR2X1_19 gnd vdd FILL
XFILL_76_DFFSR_99 gnd vdd FILL
XFILL_3_NAND2X1_53 gnd vdd FILL
XOAI21X1_8 MUX2X1_5/A OAI21X1_8/B OAI21X1_8/C gnd OAI21X1_8/Y vdd OAI21X1
XFILL_3_NAND2X1_64 gnd vdd FILL
XFILL_3_NAND2X1_75 gnd vdd FILL
XFILL_11_BUFX4_7 gnd vdd FILL
XFILL_3_NAND2X1_86 gnd vdd FILL
XFILL_45_DFFSR_10 gnd vdd FILL
XFILL_45_DFFSR_21 gnd vdd FILL
XFILL_45_DFFSR_32 gnd vdd FILL
XFILL_45_DFFSR_43 gnd vdd FILL
XFILL_16_NOR3X1_7 gnd vdd FILL
XFILL_11_CLKBUF1_17 gnd vdd FILL
XFILL_8_NOR2X1_18 gnd vdd FILL
XFILL_11_CLKBUF1_28 gnd vdd FILL
XFILL_45_DFFSR_54 gnd vdd FILL
XFILL_8_NOR2X1_29 gnd vdd FILL
XFILL_45_DFFSR_65 gnd vdd FILL
XFILL_11_CLKBUF1_39 gnd vdd FILL
XFILL_45_DFFSR_76 gnd vdd FILL
XFILL_58_5_0 gnd vdd FILL
XFILL_45_DFFSR_87 gnd vdd FILL
XFILL_45_DFFSR_98 gnd vdd FILL
XFILL_5_2_2 gnd vdd FILL
XFILL_85_DFFSR_20 gnd vdd FILL
XFILL_85_DFFSR_31 gnd vdd FILL
XFILL_85_DFFSR_42 gnd vdd FILL
XFILL_85_DFFSR_53 gnd vdd FILL
XFILL_85_DFFSR_64 gnd vdd FILL
XFILL_29_CLKBUF1_30 gnd vdd FILL
XFILL_14_DFFSR_20 gnd vdd FILL
XFILL_29_CLKBUF1_41 gnd vdd FILL
XFILL_14_DFFSR_31 gnd vdd FILL
XFILL_85_DFFSR_75 gnd vdd FILL
XFILL_85_DFFSR_86 gnd vdd FILL
XFILL_14_DFFSR_42 gnd vdd FILL
XFILL_14_DFFSR_53 gnd vdd FILL
XFILL_85_DFFSR_97 gnd vdd FILL
XFILL_14_DFFSR_64 gnd vdd FILL
XFILL_14_DFFSR_75 gnd vdd FILL
XFILL_14_DFFSR_86 gnd vdd FILL
XFILL_14_DFFSR_97 gnd vdd FILL
XFILL_30_DFFSR_204 gnd vdd FILL
XFILL_30_DFFSR_215 gnd vdd FILL
XOAI22X1_10 INVX1_212/Y OAI22X1_48/B INVX1_216/Y OAI22X1_48/D gnd NOR2X1_63/A vdd
+ OAI22X1
XFILL_7_AOI21X1_20 gnd vdd FILL
XFILL_54_DFFSR_30 gnd vdd FILL
XFILL_30_DFFSR_226 gnd vdd FILL
XOAI22X1_21 INVX1_222/Y OAI22X1_9/B INVX1_226/Y OAI22X1_9/D gnd NOR2X1_82/B vdd OAI22X1
XFILL_41_4_0 gnd vdd FILL
XFILL_30_DFFSR_237 gnd vdd FILL
XFILL_7_AOI21X1_31 gnd vdd FILL
XFILL_54_DFFSR_41 gnd vdd FILL
XOAI22X1_32 INVX1_49/Y OAI22X1_32/B INVX1_53/Y OAI22X1_32/D gnd NOR2X1_96/A vdd OAI22X1
XFILL_25_NOR3X1_5 gnd vdd FILL
XFILL_7_AOI21X1_42 gnd vdd FILL
XOAI22X1_43 INVX1_88/Y OAI22X1_8/B INVX1_84/Y OAI22X1_3/D gnd OAI22X1_43/Y vdd OAI22X1
XFILL_54_DFFSR_52 gnd vdd FILL
XFILL_54_DFFSR_63 gnd vdd FILL
XFILL_30_DFFSR_248 gnd vdd FILL
XFILL_13_1_2 gnd vdd FILL
XFILL_7_AOI21X1_53 gnd vdd FILL
XFILL_54_DFFSR_74 gnd vdd FILL
XFILL_17_OAI22X1_11 gnd vdd FILL
XFILL_30_DFFSR_259 gnd vdd FILL
XFILL_17_OAI22X1_22 gnd vdd FILL
XFILL_7_AOI21X1_64 gnd vdd FILL
XFILL_54_DFFSR_85 gnd vdd FILL
XFILL_7_AOI21X1_75 gnd vdd FILL
XFILL_17_OAI22X1_33 gnd vdd FILL
XFILL_83_DFFSR_190 gnd vdd FILL
XFILL_54_DFFSR_96 gnd vdd FILL
XFILL_17_OAI22X1_44 gnd vdd FILL
XFILL_34_DFFSR_203 gnd vdd FILL
XFILL_34_DFFSR_214 gnd vdd FILL
XFILL_34_DFFSR_225 gnd vdd FILL
XFILL_34_DFFSR_236 gnd vdd FILL
XFILL_34_DFFSR_1 gnd vdd FILL
XFILL_34_DFFSR_247 gnd vdd FILL
XFILL_3_DFFSR_260 gnd vdd FILL
XFILL_1_CLKBUF1_12 gnd vdd FILL
XFILL_3_DFFSR_271 gnd vdd FILL
XFILL_34_DFFSR_258 gnd vdd FILL
XFILL_34_DFFSR_269 gnd vdd FILL
XFILL_1_CLKBUF1_23 gnd vdd FILL
XFILL_0_MUX2X1_16 gnd vdd FILL
XFILL_23_DFFSR_40 gnd vdd FILL
XFILL_1_CLKBUF1_34 gnd vdd FILL
XFILL_0_MUX2X1_27 gnd vdd FILL
XFILL_38_DFFSR_202 gnd vdd FILL
XFILL_23_DFFSR_51 gnd vdd FILL
XFILL_61_DFFSR_103 gnd vdd FILL
XFILL_61_DFFSR_114 gnd vdd FILL
XFILL_23_DFFSR_62 gnd vdd FILL
XFILL_0_MUX2X1_38 gnd vdd FILL
XFILL_38_DFFSR_213 gnd vdd FILL
XFILL_23_DFFSR_73 gnd vdd FILL
XFILL_0_MUX2X1_49 gnd vdd FILL
XFILL_61_DFFSR_125 gnd vdd FILL
XFILL_23_DFFSR_84 gnd vdd FILL
XFILL_38_DFFSR_224 gnd vdd FILL
XFILL_61_DFFSR_136 gnd vdd FILL
XFILL_38_DFFSR_235 gnd vdd FILL
XFILL_23_DFFSR_95 gnd vdd FILL
XFILL_38_DFFSR_246 gnd vdd FILL
XFILL_61_DFFSR_147 gnd vdd FILL
XFILL_61_DFFSR_158 gnd vdd FILL
XFILL_8_NOR3X1_6 gnd vdd FILL
XFILL_38_DFFSR_257 gnd vdd FILL
XFILL_7_DFFSR_270 gnd vdd FILL
XFILL_61_DFFSR_169 gnd vdd FILL
XFILL_38_DFFSR_268 gnd vdd FILL
XFILL_4_MUX2X1_15 gnd vdd FILL
XFILL_4_MUX2X1_26 gnd vdd FILL
XFILL_65_DFFSR_102 gnd vdd FILL
XFILL_63_DFFSR_50 gnd vdd FILL
XFILL_4_MUX2X1_37 gnd vdd FILL
XFILL_65_DFFSR_113 gnd vdd FILL
XFILL_63_DFFSR_61 gnd vdd FILL
XFILL_65_DFFSR_124 gnd vdd FILL
XFILL_10_OAI21X1_13 gnd vdd FILL
XFILL_4_MUX2X1_48 gnd vdd FILL
XFILL_63_DFFSR_72 gnd vdd FILL
XFILL_63_DFFSR_83 gnd vdd FILL
XFILL_10_OAI21X1_24 gnd vdd FILL
XFILL_65_DFFSR_135 gnd vdd FILL
XFILL_4_MUX2X1_59 gnd vdd FILL
XFILL_63_DFFSR_94 gnd vdd FILL
XFILL_10_OAI21X1_35 gnd vdd FILL
XFILL_65_DFFSR_146 gnd vdd FILL
XFILL_10_OAI21X1_46 gnd vdd FILL
XFILL_65_DFFSR_157 gnd vdd FILL
XFILL_3_5 gnd vdd FILL
XFILL_65_DFFSR_168 gnd vdd FILL
XFILL_65_DFFSR_179 gnd vdd FILL
XFILL_8_MUX2X1_14 gnd vdd FILL
XFILL_8_MUX2X1_25 gnd vdd FILL
XFILL_6_DFFSR_30 gnd vdd FILL
XFILL_69_DFFSR_101 gnd vdd FILL
XFILL_49_5_0 gnd vdd FILL
XFILL_8_MUX2X1_36 gnd vdd FILL
XFILL_56_DFFSR_5 gnd vdd FILL
XFILL_6_DFFSR_41 gnd vdd FILL
XFILL_69_DFFSR_112 gnd vdd FILL
XFILL_8_MUX2X1_47 gnd vdd FILL
XFILL_6_DFFSR_52 gnd vdd FILL
XFILL_69_DFFSR_123 gnd vdd FILL
XFILL_6_DFFSR_63 gnd vdd FILL
XFILL_69_DFFSR_134 gnd vdd FILL
XFILL_8_MUX2X1_58 gnd vdd FILL
XFILL_8_MUX2X1_69 gnd vdd FILL
XFILL_6_DFFSR_74 gnd vdd FILL
XFILL_12_OAI21X1_2 gnd vdd FILL
XFILL_69_DFFSR_145 gnd vdd FILL
XFILL_6_DFFSR_85 gnd vdd FILL
XFILL_69_DFFSR_156 gnd vdd FILL
XFILL_32_DFFSR_60 gnd vdd FILL
XFILL_69_DFFSR_167 gnd vdd FILL
XFILL_6_DFFSR_96 gnd vdd FILL
XFILL_32_DFFSR_71 gnd vdd FILL
XFILL_32_DFFSR_82 gnd vdd FILL
XFILL_69_DFFSR_178 gnd vdd FILL
XFILL_32_DFFSR_93 gnd vdd FILL
XFILL_7_OAI22X1_50 gnd vdd FILL
XFILL_69_DFFSR_189 gnd vdd FILL
XFILL_45_5 gnd vdd FILL
XFILL_63_0_2 gnd vdd FILL
XFILL_0_INVX1_220 gnd vdd FILL
XFILL_38_4 gnd vdd FILL
XFILL_72_DFFSR_70 gnd vdd FILL
XFILL_72_DFFSR_81 gnd vdd FILL
XFILL_72_DFFSR_92 gnd vdd FILL
XFILL_20_MUX2X1_13 gnd vdd FILL
XFILL_20_MUX2X1_24 gnd vdd FILL
XFILL_32_4_0 gnd vdd FILL
XFILL_20_MUX2X1_35 gnd vdd FILL
XFILL_20_MUX2X1_46 gnd vdd FILL
XFILL_20_MUX2X1_57 gnd vdd FILL
XFILL_20_MUX2X1_68 gnd vdd FILL
XFILL_20_MUX2X1_79 gnd vdd FILL
XFILL_78_DFFSR_9 gnd vdd FILL
XFILL_0_OAI21X1_30 gnd vdd FILL
XFILL_50_DFFSR_190 gnd vdd FILL
XFILL_41_DFFSR_80 gnd vdd FILL
XFILL_0_OAI21X1_41 gnd vdd FILL
XFILL_41_DFFSR_91 gnd vdd FILL
XFILL_81_DFFSR_90 gnd vdd FILL
XFILL_10_DFFSR_90 gnd vdd FILL
XFILL_32_DFFSR_102 gnd vdd FILL
XFILL_32_DFFSR_113 gnd vdd FILL
XFILL_32_DFFSR_124 gnd vdd FILL
XFILL_32_DFFSR_135 gnd vdd FILL
XFILL_32_DFFSR_146 gnd vdd FILL
XFILL_32_DFFSR_157 gnd vdd FILL
XFILL_1_DFFSR_170 gnd vdd FILL
XFILL_32_DFFSR_168 gnd vdd FILL
XFILL_1_DFFSR_181 gnd vdd FILL
XFILL_32_DFFSR_179 gnd vdd FILL
XFILL_1_DFFSR_192 gnd vdd FILL
XFILL_36_DFFSR_101 gnd vdd FILL
XFILL_36_DFFSR_112 gnd vdd FILL
XFILL_2_NAND3X1_17 gnd vdd FILL
XFILL_36_DFFSR_123 gnd vdd FILL
XFILL_36_DFFSR_134 gnd vdd FILL
XFILL_2_NAND3X1_28 gnd vdd FILL
XFILL_36_DFFSR_145 gnd vdd FILL
XFILL_2_NAND3X1_39 gnd vdd FILL
XFILL_36_DFFSR_156 gnd vdd FILL
XFILL_54_0_2 gnd vdd FILL
XFILL_5_DFFSR_180 gnd vdd FILL
XFILL_36_DFFSR_167 gnd vdd FILL
XFILL_36_DFFSR_178 gnd vdd FILL
XFILL_5_DFFSR_191 gnd vdd FILL
XFILL_6_NAND2X1_19 gnd vdd FILL
XFILL_36_DFFSR_189 gnd vdd FILL
XFILL_15_BUFX4_8 gnd vdd FILL
XFILL_23_4_0 gnd vdd FILL
XFILL_9_DFFSR_190 gnd vdd FILL
XFILL_16_MUX2X1_150 gnd vdd FILL
XFILL_16_MUX2X1_161 gnd vdd FILL
XFILL_16_MUX2X1_172 gnd vdd FILL
XFILL_16_MUX2X1_183 gnd vdd FILL
XFILL_16_MUX2X1_194 gnd vdd FILL
XFILL_82_DFFSR_202 gnd vdd FILL
XFILL_82_DFFSR_213 gnd vdd FILL
XFILL_82_DFFSR_224 gnd vdd FILL
XFILL_82_DFFSR_235 gnd vdd FILL
XFILL_82_DFFSR_246 gnd vdd FILL
XFILL_82_DFFSR_257 gnd vdd FILL
XFILL_82_DFFSR_268 gnd vdd FILL
XFILL_86_DFFSR_201 gnd vdd FILL
XFILL_86_DFFSR_212 gnd vdd FILL
XFILL_86_DFFSR_223 gnd vdd FILL
XFILL_86_DFFSR_234 gnd vdd FILL
XFILL_13_AOI21X1_8 gnd vdd FILL
XFILL_86_DFFSR_245 gnd vdd FILL
XFILL_86_DFFSR_256 gnd vdd FILL
XFILL_86_DFFSR_267 gnd vdd FILL
XFILL_11_BUFX2_4 gnd vdd FILL
XFILL_2_INVX1_140 gnd vdd FILL
XFILL_2_INVX1_151 gnd vdd FILL
XFILL_2_INVX1_162 gnd vdd FILL
XFILL_2_INVX1_173 gnd vdd FILL
XFILL_2_INVX1_184 gnd vdd FILL
XFILL_2_INVX1_195 gnd vdd FILL
XFILL_21_CLKBUF1_18 gnd vdd FILL
XFILL_21_CLKBUF1_29 gnd vdd FILL
XFILL_6_5_0 gnd vdd FILL
XFILL_6_INVX1_150 gnd vdd FILL
XFILL_38_DFFSR_2 gnd vdd FILL
XFILL_6_INVX1_161 gnd vdd FILL
XFILL_0_INVX1_18 gnd vdd FILL
XFILL_6_INVX1_172 gnd vdd FILL
XFILL_6_INVX1_183 gnd vdd FILL
XFILL_6_INVX1_194 gnd vdd FILL
XFILL_0_INVX1_29 gnd vdd FILL
XFILL_45_0_2 gnd vdd FILL
XFILL_0_OAI22X1_2 gnd vdd FILL
XFILL_14_4_0 gnd vdd FILL
XFILL_2_NOR2X1_107 gnd vdd FILL
XFILL_2_NOR2X1_118 gnd vdd FILL
XFILL_2_NOR2X1_129 gnd vdd FILL
XFILL_4_OAI22X1_1 gnd vdd FILL
XFILL_22_DFFSR_8 gnd vdd FILL
XFILL_55_DFFSR_19 gnd vdd FILL
XFILL_53_DFFSR_201 gnd vdd FILL
XFILL_53_DFFSR_212 gnd vdd FILL
XFILL_53_DFFSR_223 gnd vdd FILL
XFILL_53_DFFSR_234 gnd vdd FILL
XFILL_53_DFFSR_245 gnd vdd FILL
XFILL_53_DFFSR_256 gnd vdd FILL
XFILL_53_DFFSR_267 gnd vdd FILL
XFILL_9_NAND3X1_70 gnd vdd FILL
XFILL_9_NAND3X1_81 gnd vdd FILL
XFILL_80_DFFSR_101 gnd vdd FILL
XFILL_57_DFFSR_200 gnd vdd FILL
XFILL_9_NAND3X1_92 gnd vdd FILL
XFILL_24_DFFSR_18 gnd vdd FILL
XFILL_80_DFFSR_112 gnd vdd FILL
XFILL_57_DFFSR_211 gnd vdd FILL
XFILL_15_BUFX4_50 gnd vdd FILL
XFILL_1_2 gnd vdd FILL
XFILL_80_DFFSR_123 gnd vdd FILL
XFILL_57_DFFSR_222 gnd vdd FILL
XFILL_24_DFFSR_29 gnd vdd FILL
XFILL_80_DFFSR_134 gnd vdd FILL
XFILL_57_DFFSR_233 gnd vdd FILL
XFILL_15_BUFX4_61 gnd vdd FILL
XFILL_80_DFFSR_145 gnd vdd FILL
XFILL_57_DFFSR_244 gnd vdd FILL
XFILL_15_BUFX4_72 gnd vdd FILL
XFILL_80_DFFSR_156 gnd vdd FILL
XFILL_15_BUFX4_83 gnd vdd FILL
XFILL_57_DFFSR_255 gnd vdd FILL
XFILL_80_DFFSR_167 gnd vdd FILL
XFILL_15_BUFX4_94 gnd vdd FILL
XFILL_80_DFFSR_178 gnd vdd FILL
XFILL_57_DFFSR_266 gnd vdd FILL
XFILL_12_CLKBUF1_7 gnd vdd FILL
XFILL_3_OAI21X1_18 gnd vdd FILL
XFILL_3_OAI21X1_29 gnd vdd FILL
XFILL_84_DFFSR_100 gnd vdd FILL
XFILL_80_DFFSR_189 gnd vdd FILL
XFILL_0_DFFSR_204 gnd vdd FILL
XFILL_0_DFFSR_215 gnd vdd FILL
XFILL_64_DFFSR_17 gnd vdd FILL
XFILL_84_DFFSR_111 gnd vdd FILL
XFILL_64_DFFSR_28 gnd vdd FILL
XFILL_0_DFFSR_226 gnd vdd FILL
XFILL_84_DFFSR_122 gnd vdd FILL
XFILL_84_DFFSR_133 gnd vdd FILL
XFILL_50_3 gnd vdd FILL
XFILL_0_DFFSR_237 gnd vdd FILL
XFILL_64_DFFSR_39 gnd vdd FILL
XFILL_84_DFFSR_144 gnd vdd FILL
XFILL_0_DFFSR_248 gnd vdd FILL
XFILL_64_3_0 gnd vdd FILL
XFILL_84_DFFSR_155 gnd vdd FILL
XFILL_0_DFFSR_259 gnd vdd FILL
XFILL_43_2 gnd vdd FILL
XFILL_36_0_2 gnd vdd FILL
XFILL_84_DFFSR_166 gnd vdd FILL
XFILL_84_DFFSR_177 gnd vdd FILL
XFILL_16_CLKBUF1_6 gnd vdd FILL
XFILL_84_DFFSR_188 gnd vdd FILL
XFILL_4_DFFSR_203 gnd vdd FILL
XFILL_1_NAND3X1_3 gnd vdd FILL
XFILL_2_NAND2X1_50 gnd vdd FILL
XFILL_84_DFFSR_199 gnd vdd FILL
XFILL_4_DFFSR_214 gnd vdd FILL
XFILL_4_DFFSR_225 gnd vdd FILL
XFILL_2_NAND2X1_61 gnd vdd FILL
XFILL_7_DFFSR_19 gnd vdd FILL
XFILL_2_NAND2X1_72 gnd vdd FILL
XFILL_4_DFFSR_236 gnd vdd FILL
XFILL_4_DFFSR_247 gnd vdd FILL
XFILL_2_NAND2X1_83 gnd vdd FILL
XFILL_2_NAND2X1_94 gnd vdd FILL
XFILL_12_BUFX4_101 gnd vdd FILL
XFILL_33_DFFSR_16 gnd vdd FILL
XFILL_4_DFFSR_258 gnd vdd FILL
XFILL_4_DFFSR_269 gnd vdd FILL
XFILL_33_DFFSR_27 gnd vdd FILL
XFILL_33_DFFSR_38 gnd vdd FILL
XFILL_8_DFFSR_202 gnd vdd FILL
XFILL_33_DFFSR_49 gnd vdd FILL
XFILL_10_CLKBUF1_14 gnd vdd FILL
XFILL_5_NAND3X1_2 gnd vdd FILL
XFILL_10_CLKBUF1_25 gnd vdd FILL
XFILL_8_DFFSR_213 gnd vdd FILL
XFILL_10_CLKBUF1_36 gnd vdd FILL
XFILL_8_DFFSR_224 gnd vdd FILL
XFILL_8_DFFSR_235 gnd vdd FILL
XFILL_8_DFFSR_246 gnd vdd FILL
XFILL_8_DFFSR_257 gnd vdd FILL
XFILL_73_DFFSR_15 gnd vdd FILL
XFILL_8_DFFSR_268 gnd vdd FILL
XFILL_73_DFFSR_26 gnd vdd FILL
XFILL_73_DFFSR_37 gnd vdd FILL
XFILL_73_DFFSR_48 gnd vdd FILL
XFILL_16_MUX2X1_5 gnd vdd FILL
XFILL_9_NAND3X1_1 gnd vdd FILL
XFILL_73_DFFSR_59 gnd vdd FILL
XFILL_7_BUFX4_60 gnd vdd FILL
XFILL_7_BUFX4_71 gnd vdd FILL
XFILL_42_DFFSR_14 gnd vdd FILL
XFILL_20_DFFSR_201 gnd vdd FILL
XFILL_42_DFFSR_25 gnd vdd FILL
XFILL_42_DFFSR_36 gnd vdd FILL
XFILL_20_DFFSR_212 gnd vdd FILL
XFILL_19_MUX2X1_105 gnd vdd FILL
XFILL_7_BUFX4_82 gnd vdd FILL
XFILL_10_NOR2X1_14 gnd vdd FILL
XFILL_7_BUFX4_93 gnd vdd FILL
XFILL_10_NOR2X1_25 gnd vdd FILL
XFILL_19_MUX2X1_116 gnd vdd FILL
XFILL_20_DFFSR_223 gnd vdd FILL
XFILL_42_DFFSR_47 gnd vdd FILL
XFILL_20_DFFSR_234 gnd vdd FILL
XFILL_42_DFFSR_58 gnd vdd FILL
XFILL_19_MUX2X1_127 gnd vdd FILL
XFILL_1_AOI22X1_8 gnd vdd FILL
XFILL_19_MUX2X1_138 gnd vdd FILL
XFILL_20_DFFSR_245 gnd vdd FILL
XFILL_10_NOR2X1_36 gnd vdd FILL
XFILL_10_NOR2X1_47 gnd vdd FILL
XFILL_6_AOI21X1_50 gnd vdd FILL
XFILL_42_DFFSR_69 gnd vdd FILL
XFILL_19_MUX2X1_149 gnd vdd FILL
XFILL_10_NOR2X1_58 gnd vdd FILL
XFILL_20_DFFSR_256 gnd vdd FILL
XFILL_6_AOI21X1_61 gnd vdd FILL
XFILL_20_DFFSR_267 gnd vdd FILL
XFILL_10_NOR2X1_69 gnd vdd FILL
XFILL_82_DFFSR_13 gnd vdd FILL
XFILL_6_AOI21X1_72 gnd vdd FILL
XFILL_16_OAI22X1_30 gnd vdd FILL
XFILL_16_OAI22X1_41 gnd vdd FILL
XFILL_1_INVX1_207 gnd vdd FILL
XFILL_24_DFFSR_200 gnd vdd FILL
XFILL_82_DFFSR_24 gnd vdd FILL
XFILL_1_INVX1_218 gnd vdd FILL
XFILL_24_DFFSR_211 gnd vdd FILL
XFILL_82_DFFSR_35 gnd vdd FILL
XFILL_24_DFFSR_222 gnd vdd FILL
XFILL_82_DFFSR_46 gnd vdd FILL
XFILL_11_DFFSR_13 gnd vdd FILL
XFILL_82_DFFSR_57 gnd vdd FILL
XFILL_24_DFFSR_233 gnd vdd FILL
XFILL_5_AOI22X1_7 gnd vdd FILL
XFILL_82_DFFSR_68 gnd vdd FILL
XFILL_24_DFFSR_244 gnd vdd FILL
XFILL_7_DFFSR_1 gnd vdd FILL
XFILL_11_DFFSR_24 gnd vdd FILL
XFILL_24_DFFSR_255 gnd vdd FILL
XFILL_11_DFFSR_35 gnd vdd FILL
XFILL_82_DFFSR_79 gnd vdd FILL
XFILL_9_NOR2X1_160 gnd vdd FILL
XFILL_0_CLKBUF1_20 gnd vdd FILL
XFILL_11_DFFSR_46 gnd vdd FILL
XFILL_24_DFFSR_266 gnd vdd FILL
XFILL_11_DFFSR_57 gnd vdd FILL
XFILL_0_CLKBUF1_31 gnd vdd FILL
XFILL_9_NOR2X1_171 gnd vdd FILL
XFILL_5_INVX1_206 gnd vdd FILL
XFILL_11_DFFSR_68 gnd vdd FILL
XFILL_51_DFFSR_100 gnd vdd FILL
XFILL_0_CLKBUF1_42 gnd vdd FILL
XFILL_9_NOR2X1_182 gnd vdd FILL
XFILL_9_NOR2X1_6 gnd vdd FILL
XFILL_55_3_0 gnd vdd FILL
XFILL_28_DFFSR_210 gnd vdd FILL
XFILL_9_NOR2X1_193 gnd vdd FILL
XFILL_51_DFFSR_111 gnd vdd FILL
XFILL_5_INVX1_217 gnd vdd FILL
XFILL_11_DFFSR_79 gnd vdd FILL
XFILL_5_INVX1_228 gnd vdd FILL
XFILL_51_DFFSR_122 gnd vdd FILL
XFILL_27_0_2 gnd vdd FILL
XFILL_9_AOI22X1_6 gnd vdd FILL
XFILL_51_DFFSR_133 gnd vdd FILL
XFILL_2_0_2 gnd vdd FILL
XFILL_28_DFFSR_221 gnd vdd FILL
XFILL_51_DFFSR_12 gnd vdd FILL
XFILL_28_DFFSR_232 gnd vdd FILL
XFILL_28_DFFSR_243 gnd vdd FILL
XFILL_51_DFFSR_144 gnd vdd FILL
XFILL_51_DFFSR_23 gnd vdd FILL
XFILL_51_DFFSR_155 gnd vdd FILL
XFILL_28_DFFSR_254 gnd vdd FILL
XFILL_51_DFFSR_34 gnd vdd FILL
XFILL_51_DFFSR_166 gnd vdd FILL
XFILL_2_BUFX2_7 gnd vdd FILL
XFILL_51_DFFSR_177 gnd vdd FILL
XFILL_22_NOR3X1_9 gnd vdd FILL
XFILL_51_DFFSR_45 gnd vdd FILL
XFILL_28_DFFSR_265 gnd vdd FILL
XFILL_51_DFFSR_56 gnd vdd FILL
XFILL_51_DFFSR_67 gnd vdd FILL
XFILL_51_DFFSR_188 gnd vdd FILL
XFILL_51_DFFSR_78 gnd vdd FILL
XFILL_55_DFFSR_110 gnd vdd FILL
XFILL_51_DFFSR_199 gnd vdd FILL
XFILL_55_DFFSR_121 gnd vdd FILL
XFILL_51_DFFSR_89 gnd vdd FILL
XFILL_55_DFFSR_132 gnd vdd FILL
XFILL_55_DFFSR_143 gnd vdd FILL
XFILL_55_DFFSR_154 gnd vdd FILL
XFILL_8_MUX2X1_4 gnd vdd FILL
XFILL_55_DFFSR_165 gnd vdd FILL
XFILL_55_DFFSR_176 gnd vdd FILL
XFILL_9_MUX2X1_100 gnd vdd FILL
XFILL_20_DFFSR_11 gnd vdd FILL
XFILL_55_DFFSR_187 gnd vdd FILL
XFILL_9_MUX2X1_111 gnd vdd FILL
XFILL_61_DFFSR_6 gnd vdd FILL
XFILL_20_DFFSR_22 gnd vdd FILL
XFILL_55_DFFSR_198 gnd vdd FILL
XFILL_20_DFFSR_33 gnd vdd FILL
XFILL_9_MUX2X1_122 gnd vdd FILL
XFILL_59_DFFSR_120 gnd vdd FILL
XFILL_59_DFFSR_131 gnd vdd FILL
XFILL_9_MUX2X1_133 gnd vdd FILL
XFILL_20_DFFSR_44 gnd vdd FILL
XFILL_9_MUX2X1_144 gnd vdd FILL
XFILL_20_DFFSR_55 gnd vdd FILL
XFILL_59_DFFSR_142 gnd vdd FILL
XFILL_9_MUX2X1_155 gnd vdd FILL
XFILL_20_DFFSR_66 gnd vdd FILL
XFILL_20_DFFSR_77 gnd vdd FILL
XFILL_59_DFFSR_153 gnd vdd FILL
XFILL_13_OR2X2_1 gnd vdd FILL
XFILL_20_DFFSR_88 gnd vdd FILL
XFILL_9_MUX2X1_166 gnd vdd FILL
XFILL_59_DFFSR_164 gnd vdd FILL
XFILL_59_DFFSR_175 gnd vdd FILL
XFILL_9_MUX2X1_177 gnd vdd FILL
XFILL_2_DFFSR_102 gnd vdd FILL
XFILL_20_DFFSR_99 gnd vdd FILL
XFILL_59_DFFSR_186 gnd vdd FILL
XFILL_9_MUX2X1_188 gnd vdd FILL
XFILL_60_DFFSR_10 gnd vdd FILL
XFILL_60_DFFSR_21 gnd vdd FILL
XFILL_59_DFFSR_197 gnd vdd FILL
XFILL_2_DFFSR_113 gnd vdd FILL
XFILL_2_DFFSR_124 gnd vdd FILL
XFILL_60_DFFSR_32 gnd vdd FILL
XFILL_60_DFFSR_43 gnd vdd FILL
XFILL_2_DFFSR_135 gnd vdd FILL
XFILL_31_NOR3X1_7 gnd vdd FILL
XFILL_2_DFFSR_146 gnd vdd FILL
XFILL_60_DFFSR_54 gnd vdd FILL
XFILL_2_DFFSR_157 gnd vdd FILL
XFILL_60_DFFSR_65 gnd vdd FILL
XFILL_60_DFFSR_76 gnd vdd FILL
XFILL_2_DFFSR_168 gnd vdd FILL
XDFFSR_90 DFFSR_90/Q DFFSR_90/CLK DFFSR_90/R vdd DFFSR_90/D gnd vdd DFFSR
XFILL_2_DFFSR_179 gnd vdd FILL
XFILL_60_DFFSR_87 gnd vdd FILL
XFILL_60_DFFSR_98 gnd vdd FILL
XFILL_6_DFFSR_101 gnd vdd FILL
XFILL_10_MUX2X1_10 gnd vdd FILL
XFILL_6_DFFSR_112 gnd vdd FILL
XFILL_10_MUX2X1_21 gnd vdd FILL
XFILL_3_DFFSR_12 gnd vdd FILL
XFILL_6_DFFSR_123 gnd vdd FILL
XFILL_6_DFFSR_134 gnd vdd FILL
XFILL_10_MUX2X1_32 gnd vdd FILL
XFILL_3_DFFSR_23 gnd vdd FILL
XFILL_1_BUFX4_1 gnd vdd FILL
XFILL_3_DFFSR_34 gnd vdd FILL
XFILL_6_DFFSR_145 gnd vdd FILL
XFILL_10_MUX2X1_43 gnd vdd FILL
XFILL_6_DFFSR_156 gnd vdd FILL
XFILL_26_DFFSR_9 gnd vdd FILL
XFILL_10_MUX2X1_54 gnd vdd FILL
XFILL_3_DFFSR_45 gnd vdd FILL
XFILL_11_NAND3X1_19 gnd vdd FILL
XFILL_3_DFFSR_56 gnd vdd FILL
XFILL_6_DFFSR_167 gnd vdd FILL
XFILL_10_MUX2X1_65 gnd vdd FILL
XFILL_6_DFFSR_178 gnd vdd FILL
XFILL_10_MUX2X1_76 gnd vdd FILL
XFILL_3_DFFSR_67 gnd vdd FILL
XFILL_10_MUX2X1_87 gnd vdd FILL
XFILL_3_DFFSR_78 gnd vdd FILL
XFILL_6_DFFSR_189 gnd vdd FILL
XFILL_3_DFFSR_89 gnd vdd FILL
XFILL_10_MUX2X1_98 gnd vdd FILL
XFILL_14_MUX2X1_20 gnd vdd FILL
XFILL_31_CLKBUF1_19 gnd vdd FILL
XFILL_14_MUX2X1_31 gnd vdd FILL
XFILL_14_MUX2X1_42 gnd vdd FILL
XFILL_14_MUX2X1_53 gnd vdd FILL
XFILL_14_MUX2X1_64 gnd vdd FILL
XFILL_2_NOR3X1_13 gnd vdd FILL
XFILL_14_MUX2X1_75 gnd vdd FILL
XFILL_46_3_0 gnd vdd FILL
XFILL_14_MUX2X1_86 gnd vdd FILL
XFILL_18_0_2 gnd vdd FILL
XFILL_2_NOR3X1_24 gnd vdd FILL
XFILL_14_MUX2X1_97 gnd vdd FILL
XFILL_2_NOR3X1_35 gnd vdd FILL
XFILL_2_NOR3X1_46 gnd vdd FILL
XFILL_18_MUX2X1_30 gnd vdd FILL
XFILL_18_MUX2X1_41 gnd vdd FILL
XFILL_18_MUX2X1_52 gnd vdd FILL
XFILL_0_INVX1_5 gnd vdd FILL
XFILL_18_MUX2X1_63 gnd vdd FILL
XFILL_6_NOR3X1_12 gnd vdd FILL
XFILL_18_MUX2X1_74 gnd vdd FILL
XFILL_18_MUX2X1_85 gnd vdd FILL
XFILL_18_MUX2X1_96 gnd vdd FILL
XFILL_6_NOR3X1_23 gnd vdd FILL
XFILL_22_7 gnd vdd FILL
XFILL_6_NOR3X1_34 gnd vdd FILL
XFILL_6_NOR3X1_45 gnd vdd FILL
XFILL_22_DFFSR_110 gnd vdd FILL
XFILL_22_DFFSR_121 gnd vdd FILL
XFILL_22_DFFSR_132 gnd vdd FILL
XFILL_30_7_1 gnd vdd FILL
XFILL_22_DFFSR_143 gnd vdd FILL
XFILL_22_DFFSR_154 gnd vdd FILL
XFILL_22_DFFSR_165 gnd vdd FILL
XFILL_22_DFFSR_176 gnd vdd FILL
XFILL_3_INVX1_105 gnd vdd FILL
XFILL_22_DFFSR_187 gnd vdd FILL
XFILL_3_INVX1_116 gnd vdd FILL
XFILL_3_INVX1_127 gnd vdd FILL
XFILL_22_DFFSR_198 gnd vdd FILL
XFILL_26_DFFSR_120 gnd vdd FILL
XFILL_1_NAND3X1_14 gnd vdd FILL
XFILL_26_DFFSR_131 gnd vdd FILL
XFILL_1_NAND3X1_25 gnd vdd FILL
XFILL_3_INVX1_138 gnd vdd FILL
XFILL_26_DFFSR_142 gnd vdd FILL
XFILL_3_INVX1_149 gnd vdd FILL
XFILL_1_NAND3X1_36 gnd vdd FILL
XFILL_26_DFFSR_153 gnd vdd FILL
XFILL_1_NAND3X1_47 gnd vdd FILL
XFILL_1_INVX4_1 gnd vdd FILL
XFILL_1_NAND3X1_58 gnd vdd FILL
XFILL_26_DFFSR_164 gnd vdd FILL
XFILL_1_NAND3X1_69 gnd vdd FILL
XFILL_26_DFFSR_175 gnd vdd FILL
XFILL_5_NAND2X1_16 gnd vdd FILL
XFILL_7_INVX1_104 gnd vdd FILL
XFILL_5_NAND2X1_27 gnd vdd FILL
XFILL_26_DFFSR_186 gnd vdd FILL
XFILL_7_INVX1_115 gnd vdd FILL
XFILL_5_NAND2X1_38 gnd vdd FILL
XFILL_5_NAND2X1_49 gnd vdd FILL
XFILL_7_INVX1_126 gnd vdd FILL
XFILL_26_DFFSR_197 gnd vdd FILL
XINVX1_140 BUFX2_9/A gnd INVX1_140/Y vdd INVX1
XINVX1_151 INVX1_151/A gnd NOR2X1_62/A vdd INVX1
XFILL_7_INVX1_137 gnd vdd FILL
XINVX1_162 INVX1_162/A gnd INVX1_162/Y vdd INVX1
XFILL_7_INVX1_148 gnd vdd FILL
XFILL_7_INVX1_159 gnd vdd FILL
XINVX1_173 INVX1_173/A gnd INVX1_173/Y vdd INVX1
XINVX1_184 INVX1_184/A gnd INVX1_184/Y vdd INVX1
XINVX1_195 DFFSR_97/Q gnd INVX1_195/Y vdd INVX1
XFILL_22_NOR3X1_10 gnd vdd FILL
XFILL_22_NOR3X1_21 gnd vdd FILL
XFILL_22_NOR3X1_32 gnd vdd FILL
XFILL_15_MUX2X1_180 gnd vdd FILL
XFILL_22_NOR3X1_43 gnd vdd FILL
XFILL_15_MUX2X1_191 gnd vdd FILL
XFILL_72_DFFSR_210 gnd vdd FILL
XFILL_72_DFFSR_221 gnd vdd FILL
XFILL_72_DFFSR_232 gnd vdd FILL
XFILL_72_DFFSR_243 gnd vdd FILL
XFILL_72_DFFSR_254 gnd vdd FILL
XFILL_26_NOR3X1_20 gnd vdd FILL
XFILL_72_DFFSR_265 gnd vdd FILL
XFILL_26_NOR3X1_31 gnd vdd FILL
XFILL_26_NOR3X1_42 gnd vdd FILL
XFILL_37_3_0 gnd vdd FILL
XFILL_76_DFFSR_220 gnd vdd FILL
XFILL_11_NOR2X1_109 gnd vdd FILL
XFILL_76_DFFSR_231 gnd vdd FILL
XFILL_1_NOR3X1_3 gnd vdd FILL
XFILL_76_DFFSR_242 gnd vdd FILL
XFILL_76_DFFSR_253 gnd vdd FILL
XFILL_76_DFFSR_264 gnd vdd FILL
XFILL_31_CLKBUF1_5 gnd vdd FILL
XFILL_76_DFFSR_275 gnd vdd FILL
XFILL_9_AOI21X1_16 gnd vdd FILL
XFILL_9_OAI22X1_9 gnd vdd FILL
XFILL_9_AOI21X1_27 gnd vdd FILL
XFILL_9_AOI21X1_38 gnd vdd FILL
XFILL_9_AOI21X1_49 gnd vdd FILL
XFILL_19_OAI22X1_18 gnd vdd FILL
XFILL_35_CLKBUF1_4 gnd vdd FILL
XFILL_21_7_1 gnd vdd FILL
XFILL_19_OAI22X1_29 gnd vdd FILL
XFILL_20_CLKBUF1_15 gnd vdd FILL
XFILL_20_CLKBUF1_26 gnd vdd FILL
XFILL_20_2_0 gnd vdd FILL
XFILL_20_CLKBUF1_37 gnd vdd FILL
XFILL_43_DFFSR_3 gnd vdd FILL
XFILL_3_CLKBUF1_19 gnd vdd FILL
XFILL_58_DFFSR_209 gnd vdd FILL
XFILL_6_BUFX2_8 gnd vdd FILL
XFILL_85_DFFSR_109 gnd vdd FILL
XFILL_1_NOR2X1_104 gnd vdd FILL
XFILL_1_NOR2X1_115 gnd vdd FILL
XFILL_1_NOR2X1_126 gnd vdd FILL
XFILL_1_NOR2X1_137 gnd vdd FILL
XFILL_1_NOR2X1_148 gnd vdd FILL
XFILL_1_NOR2X1_159 gnd vdd FILL
XFILL_65_DFFSR_7 gnd vdd FILL
XFILL_8_BUFX4_16 gnd vdd FILL
XFILL_11_NAND2X1_30 gnd vdd FILL
XFILL_8_BUFX4_27 gnd vdd FILL
XFILL_11_NAND2X1_41 gnd vdd FILL
XFILL_8_BUFX4_38 gnd vdd FILL
XFILL_11_NAND2X1_52 gnd vdd FILL
XFILL_8_BUFX4_49 gnd vdd FILL
XFILL_11_NAND2X1_63 gnd vdd FILL
XFILL_9_OAI22X1_13 gnd vdd FILL
XFILL_11_NAND2X1_74 gnd vdd FILL
XFILL_11_NAND2X1_85 gnd vdd FILL
XFILL_9_OAI22X1_24 gnd vdd FILL
XFILL_28_3_0 gnd vdd FILL
XFILL_9_OAI22X1_35 gnd vdd FILL
XFILL_3_3_0 gnd vdd FILL
XFILL_11_NAND2X1_96 gnd vdd FILL
XFILL_9_OAI22X1_46 gnd vdd FILL
XFILL_43_DFFSR_220 gnd vdd FILL
XFILL_43_DFFSR_231 gnd vdd FILL
XFILL_43_DFFSR_242 gnd vdd FILL
XFILL_43_DFFSR_253 gnd vdd FILL
XFILL_43_DFFSR_264 gnd vdd FILL
XNAND3X1_104 INVX1_107/A BUFX4_58/Y AND2X2_6/Y gnd NAND3X1_106/B vdd NAND3X1
XFILL_43_DFFSR_275 gnd vdd FILL
XFILL_2_NOR2X1_90 gnd vdd FILL
XNAND3X1_115 NOR2X1_46/A BUFX4_91/Y NOR2X1_38/Y gnd NAND3X1_118/B vdd NAND3X1
XNAND3X1_126 NAND3X1_126/A INVX1_128/Y NOR2X1_85/Y gnd NOR2X1_91/A vdd NAND3X1
XFILL_5_BUFX4_2 gnd vdd FILL
XFILL_6_NOR2X1_204 gnd vdd FILL
XFILL_70_DFFSR_120 gnd vdd FILL
XFILL_70_DFFSR_131 gnd vdd FILL
XFILL_12_7_1 gnd vdd FILL
XFILL_47_DFFSR_230 gnd vdd FILL
XFILL_70_DFFSR_142 gnd vdd FILL
XFILL_47_DFFSR_241 gnd vdd FILL
XFILL_70_DFFSR_153 gnd vdd FILL
XFILL_11_2_0 gnd vdd FILL
XFILL_47_DFFSR_252 gnd vdd FILL
XFILL_15_AND2X2_4 gnd vdd FILL
XFILL_47_DFFSR_263 gnd vdd FILL
XFILL_70_DFFSR_164 gnd vdd FILL
XFILL_70_DFFSR_175 gnd vdd FILL
XFILL_47_DFFSR_274 gnd vdd FILL
XFILL_2_OAI21X1_15 gnd vdd FILL
XFILL_70_DFFSR_186 gnd vdd FILL
XFILL_2_OAI21X1_26 gnd vdd FILL
XFILL_70_DFFSR_197 gnd vdd FILL
XFILL_2_OAI21X1_37 gnd vdd FILL
XFILL_74_DFFSR_130 gnd vdd FILL
XFILL_2_OAI21X1_48 gnd vdd FILL
XFILL_74_DFFSR_141 gnd vdd FILL
XFILL_74_DFFSR_152 gnd vdd FILL
XFILL_15_AOI21X1_30 gnd vdd FILL
XFILL_74_DFFSR_163 gnd vdd FILL
XFILL_74_DFFSR_174 gnd vdd FILL
XFILL_15_AOI21X1_41 gnd vdd FILL
XFILL_74_DFFSR_185 gnd vdd FILL
XFILL_15_AOI21X1_52 gnd vdd FILL
XFILL_74_DFFSR_196 gnd vdd FILL
XFILL_12_BUFX4_10 gnd vdd FILL
XFILL_15_AOI21X1_63 gnd vdd FILL
XFILL_15_AOI21X1_74 gnd vdd FILL
XFILL_25_DFFSR_209 gnd vdd FILL
XFILL_12_BUFX4_21 gnd vdd FILL
XFILL_78_DFFSR_140 gnd vdd FILL
XFILL_1_NAND2X1_80 gnd vdd FILL
XFILL_4_INVX1_6 gnd vdd FILL
XFILL_12_BUFX4_32 gnd vdd FILL
XFILL_12_BUFX4_43 gnd vdd FILL
XFILL_78_DFFSR_151 gnd vdd FILL
XFILL_1_NAND2X1_91 gnd vdd FILL
XFILL_12_BUFX4_54 gnd vdd FILL
XFILL_78_DFFSR_162 gnd vdd FILL
XFILL_12_BUFX4_65 gnd vdd FILL
XFILL_78_DFFSR_173 gnd vdd FILL
XFILL_78_DFFSR_184 gnd vdd FILL
XFILL_12_BUFX4_76 gnd vdd FILL
XFILL_78_DFFSR_195 gnd vdd FILL
XFILL_12_BUFX4_87 gnd vdd FILL
XFILL_52_DFFSR_109 gnd vdd FILL
XFILL_29_DFFSR_208 gnd vdd FILL
XFILL_12_BUFX4_98 gnd vdd FILL
XFILL_29_DFFSR_219 gnd vdd FILL
XFILL_2_NAND2X1_1 gnd vdd FILL
XFILL_56_DFFSR_108 gnd vdd FILL
XFILL_56_DFFSR_119 gnd vdd FILL
XFILL_19_3_0 gnd vdd FILL
XFILL_62_6_1 gnd vdd FILL
XFILL_6_INVX1_11 gnd vdd FILL
XFILL_6_INVX1_22 gnd vdd FILL
XFILL_61_1_0 gnd vdd FILL
XFILL_6_INVX1_33 gnd vdd FILL
XFILL_18_MUX2X1_102 gnd vdd FILL
XFILL_18_MUX2X1_113 gnd vdd FILL
XFILL_10_DFFSR_220 gnd vdd FILL
XFILL_6_INVX1_44 gnd vdd FILL
XFILL_7_AND2X2_3 gnd vdd FILL
XFILL_18_MUX2X1_124 gnd vdd FILL
XFILL_6_INVX1_55 gnd vdd FILL
XFILL_10_DFFSR_231 gnd vdd FILL
XFILL_6_INVX1_66 gnd vdd FILL
XFILL_10_DFFSR_242 gnd vdd FILL
XFILL_18_MUX2X1_135 gnd vdd FILL
XFILL_20_4 gnd vdd FILL
XFILL_18_MUX2X1_146 gnd vdd FILL
XFILL_6_INVX1_77 gnd vdd FILL
XFILL_10_DFFSR_253 gnd vdd FILL
XFILL_6_INVX1_88 gnd vdd FILL
XFILL_10_DFFSR_264 gnd vdd FILL
XFILL_18_MUX2X1_157 gnd vdd FILL
XFILL_10_DFFSR_275 gnd vdd FILL
XFILL_70_DFFSR_19 gnd vdd FILL
XFILL_6_INVX1_99 gnd vdd FILL
XFILL_13_3 gnd vdd FILL
XFILL_18_MUX2X1_168 gnd vdd FILL
XFILL_5_AOI21X1_80 gnd vdd FILL
XFILL_18_MUX2X1_179 gnd vdd FILL
XFILL_13_MUX2X1_9 gnd vdd FILL
XFILL_14_DFFSR_230 gnd vdd FILL
XFILL_14_DFFSR_241 gnd vdd FILL
XDFFSR_102 DFFSR_102/Q DFFSR_94/CLK DFFSR_99/R vdd DFFSR_102/D gnd vdd DFFSR
XFILL_14_DFFSR_252 gnd vdd FILL
XFILL_4_BUFX4_20 gnd vdd FILL
XFILL_82_DFFSR_1 gnd vdd FILL
XDFFSR_113 INVX1_106/A CLKBUF1_4/Y DFFSR_90/R vdd MUX2X1_93/Y gnd vdd DFFSR
XFILL_14_DFFSR_263 gnd vdd FILL
XDFFSR_124 INVX1_107/A CLKBUF1_4/Y DFFSR_49/R vdd MUX2X1_94/Y gnd vdd DFFSR
XFILL_14_DFFSR_274 gnd vdd FILL
XFILL_4_BUFX4_31 gnd vdd FILL
XDFFSR_135 INVX1_108/A DFFSR_90/CLK BUFX4_32/Y vdd MUX2X1_95/Y gnd vdd DFFSR
XFILL_11_MUX2X1_19 gnd vdd FILL
XDFFSR_146 INVX1_100/A DFFSR_45/CLK BUFX4_13/Y vdd MUX2X1_87/Y gnd vdd DFFSR
XFILL_4_BUFX4_42 gnd vdd FILL
XFILL_8_NOR2X1_190 gnd vdd FILL
XDFFSR_157 INVX1_102/A CLKBUF1_4/Y DFFSR_90/R vdd MUX2X1_88/Y gnd vdd DFFSR
XFILL_4_BUFX4_53 gnd vdd FILL
XFILL_41_DFFSR_130 gnd vdd FILL
XFILL_4_BUFX4_64 gnd vdd FILL
XBUFX4_9 clk gnd BUFX4_9/Y vdd BUFX4
XFILL_2_AOI21X1_6 gnd vdd FILL
XDFFSR_168 INVX1_103/A DFFSR_79/CLK DFFSR_79/R vdd MUX2X1_89/Y gnd vdd DFFSR
XFILL_4_BUFX4_75 gnd vdd FILL
XDFFSR_179 INVX1_104/A CLKBUF1_7/Y BUFX4_13/Y vdd MUX2X1_91/Y gnd vdd DFFSR
XFILL_18_DFFSR_240 gnd vdd FILL
XFILL_41_DFFSR_141 gnd vdd FILL
XFILL_41_DFFSR_152 gnd vdd FILL
XFILL_18_DFFSR_251 gnd vdd FILL
XFILL_4_BUFX4_86 gnd vdd FILL
XFILL_4_BUFX4_97 gnd vdd FILL
XFILL_18_DFFSR_262 gnd vdd FILL
XFILL_41_DFFSR_163 gnd vdd FILL
XFILL_41_DFFSR_174 gnd vdd FILL
XFILL_18_DFFSR_273 gnd vdd FILL
XFILL_41_DFFSR_185 gnd vdd FILL
XFILL_15_MUX2X1_18 gnd vdd FILL
XFILL_15_MUX2X1_29 gnd vdd FILL
XFILL_41_DFFSR_196 gnd vdd FILL
XFILL_6_AOI21X1_5 gnd vdd FILL
XFILL_45_DFFSR_140 gnd vdd FILL
XFILL_45_DFFSR_151 gnd vdd FILL
XFILL_45_DFFSR_162 gnd vdd FILL
XFILL_45_DFFSR_173 gnd vdd FILL
XFILL_22_MUX2X1_7 gnd vdd FILL
XFILL_45_DFFSR_184 gnd vdd FILL
XFILL_45_DFFSR_195 gnd vdd FILL
XFILL_19_MUX2X1_17 gnd vdd FILL
XFILL_19_MUX2X1_28 gnd vdd FILL
XFILL_19_MUX2X1_39 gnd vdd FILL
XFILL_47_DFFSR_4 gnd vdd FILL
XFILL_8_MUX2X1_130 gnd vdd FILL
XFILL_8_MUX2X1_141 gnd vdd FILL
XNOR3X1_13 NOR3X1_13/A OAI22X1_7/Y OAI22X1_8/Y gnd NOR3X1_13/Y vdd NOR3X1
XFILL_49_DFFSR_150 gnd vdd FILL
XFILL_11_AOI22X1_2 gnd vdd FILL
XFILL_8_MUX2X1_152 gnd vdd FILL
XFILL_8_MUX2X1_163 gnd vdd FILL
XNOR3X1_24 NOR3X1_24/A NOR3X1_24/B NOR3X1_24/C gnd NOR3X1_24/Y vdd NOR3X1
XFILL_49_DFFSR_161 gnd vdd FILL
XNOR3X1_35 NOR3X1_35/A NOR3X1_35/B NOR3X1_35/C gnd NOR3X1_35/Y vdd NOR3X1
XFILL_49_DFFSR_172 gnd vdd FILL
XFILL_8_MUX2X1_174 gnd vdd FILL
XFILL_8_MUX2X1_185 gnd vdd FILL
XNOR3X1_46 NOR3X1_46/A NOR3X1_46/B NOR3X1_46/C gnd NOR3X1_47/A vdd NOR3X1
XFILL_49_DFFSR_183 gnd vdd FILL
XFILL_49_DFFSR_194 gnd vdd FILL
XFILL_23_DFFSR_108 gnd vdd FILL
XFILL_23_DFFSR_119 gnd vdd FILL
XFILL_53_6_1 gnd vdd FILL
XFILL_15_AOI22X1_1 gnd vdd FILL
XFILL_52_1_0 gnd vdd FILL
XFILL_5_MUX2X1_8 gnd vdd FILL
XFILL_27_DFFSR_107 gnd vdd FILL
XFILL_27_DFFSR_118 gnd vdd FILL
XFILL_27_DFFSR_129 gnd vdd FILL
XFILL_10_NAND3X1_16 gnd vdd FILL
XFILL_10_NAND3X1_27 gnd vdd FILL
XFILL_10_NAND3X1_38 gnd vdd FILL
XFILL_10_NAND3X1_49 gnd vdd FILL
XFILL_69_DFFSR_8 gnd vdd FILL
XFILL_30_CLKBUF1_16 gnd vdd FILL
XFILL_39_DFFSR_20 gnd vdd FILL
XFILL_39_DFFSR_31 gnd vdd FILL
XFILL_30_CLKBUF1_27 gnd vdd FILL
XFILL_30_CLKBUF1_38 gnd vdd FILL
XFILL_39_DFFSR_42 gnd vdd FILL
XFILL_39_DFFSR_53 gnd vdd FILL
XFILL_39_DFFSR_64 gnd vdd FILL
XFILL_39_DFFSR_75 gnd vdd FILL
XFILL_39_DFFSR_86 gnd vdd FILL
XFILL_23_NOR3X1_19 gnd vdd FILL
XFILL_39_DFFSR_97 gnd vdd FILL
XFILL_73_DFFSR_208 gnd vdd FILL
XFILL_79_DFFSR_30 gnd vdd FILL
XFILL_79_DFFSR_41 gnd vdd FILL
XFILL_73_DFFSR_219 gnd vdd FILL
XFILL_0_DFFSR_16 gnd vdd FILL
XFILL_79_DFFSR_52 gnd vdd FILL
XFILL_79_DFFSR_63 gnd vdd FILL
XFILL_0_DFFSR_27 gnd vdd FILL
XFILL_0_DFFSR_38 gnd vdd FILL
XFILL_10_NOR2X1_4 gnd vdd FILL
XFILL_79_DFFSR_74 gnd vdd FILL
XFILL_27_NOR3X1_18 gnd vdd FILL
XFILL_79_DFFSR_85 gnd vdd FILL
XFILL_0_DFFSR_49 gnd vdd FILL
XFILL_79_DFFSR_96 gnd vdd FILL
XFILL_27_NOR3X1_29 gnd vdd FILL
XFILL_77_DFFSR_207 gnd vdd FILL
XFILL_9_BUFX4_3 gnd vdd FILL
XFILL_12_DFFSR_140 gnd vdd FILL
XFILL_2_INVX1_70 gnd vdd FILL
XFILL_77_DFFSR_218 gnd vdd FILL
XFILL_77_DFFSR_229 gnd vdd FILL
XFILL_2_INVX1_81 gnd vdd FILL
XFILL_2_INVX1_92 gnd vdd FILL
XFILL_12_DFFSR_151 gnd vdd FILL
XFILL_12_DFFSR_162 gnd vdd FILL
XFILL_48_DFFSR_40 gnd vdd FILL
XFILL_12_DFFSR_173 gnd vdd FILL
XFILL_1_CLKBUF1_5 gnd vdd FILL
XFILL_19_NOR3X1_4 gnd vdd FILL
XFILL_12_DFFSR_184 gnd vdd FILL
XFILL_48_DFFSR_51 gnd vdd FILL
XFILL_48_DFFSR_62 gnd vdd FILL
XFILL_48_DFFSR_73 gnd vdd FILL
XFILL_12_DFFSR_195 gnd vdd FILL
XFILL_0_NAND3X1_11 gnd vdd FILL
XFILL_48_DFFSR_84 gnd vdd FILL
XFILL_0_NAND3X1_22 gnd vdd FILL
XFILL_48_DFFSR_95 gnd vdd FILL
XFILL_0_NAND3X1_33 gnd vdd FILL
XFILL_16_DFFSR_150 gnd vdd FILL
XFILL_0_NAND3X1_44 gnd vdd FILL
XFILL_16_DFFSR_161 gnd vdd FILL
XFILL_0_NAND3X1_55 gnd vdd FILL
XFILL_4_NAND2X1_13 gnd vdd FILL
XFILL_0_NAND3X1_66 gnd vdd FILL
XFILL_16_DFFSR_172 gnd vdd FILL
XFILL_5_CLKBUF1_4 gnd vdd FILL
XFILL_0_NAND3X1_77 gnd vdd FILL
XFILL_16_DFFSR_183 gnd vdd FILL
XFILL_4_NAND2X1_24 gnd vdd FILL
XFILL_44_6_1 gnd vdd FILL
XFILL_16_DFFSR_194 gnd vdd FILL
XFILL_4_NAND2X1_35 gnd vdd FILL
XFILL_0_NAND3X1_88 gnd vdd FILL
XFILL_4_NAND2X1_46 gnd vdd FILL
XFILL_0_NAND3X1_99 gnd vdd FILL
XFILL_4_NAND2X1_57 gnd vdd FILL
XFILL_43_1_0 gnd vdd FILL
XFILL_0_BUFX4_90 gnd vdd FILL
XFILL_4_NAND2X1_68 gnd vdd FILL
XFILL_17_DFFSR_50 gnd vdd FILL
XFILL_4_NAND2X1_79 gnd vdd FILL
XFILL_17_DFFSR_61 gnd vdd FILL
XFILL_17_DFFSR_72 gnd vdd FILL
XFILL_17_DFFSR_83 gnd vdd FILL
XFILL_9_CLKBUF1_3 gnd vdd FILL
XFILL_17_DFFSR_94 gnd vdd FILL
XFILL_28_NOR3X1_2 gnd vdd FILL
XFILL_12_NOR3X1_40 gnd vdd FILL
XFILL_12_NOR3X1_51 gnd vdd FILL
XFILL_57_DFFSR_60 gnd vdd FILL
XFILL_57_DFFSR_71 gnd vdd FILL
XFILL_57_DFFSR_82 gnd vdd FILL
XFILL_62_DFFSR_240 gnd vdd FILL
XFILL_57_DFFSR_93 gnd vdd FILL
XFILL_62_DFFSR_251 gnd vdd FILL
XFILL_62_DFFSR_262 gnd vdd FILL
XFILL_62_DFFSR_273 gnd vdd FILL
XFILL_2_NOR2X1_3 gnd vdd FILL
XFILL_16_NOR3X1_50 gnd vdd FILL
XFILL_10_NOR2X1_106 gnd vdd FILL
XFILL_10_NOR2X1_117 gnd vdd FILL
XFILL_10_NOR2X1_128 gnd vdd FILL
XFILL_66_DFFSR_250 gnd vdd FILL
XFILL_4_AOI22X1_11 gnd vdd FILL
XFILL_10_NOR2X1_139 gnd vdd FILL
XFILL_66_DFFSR_261 gnd vdd FILL
XFILL_66_DFFSR_272 gnd vdd FILL
XFILL_21_CLKBUF1_2 gnd vdd FILL
XFILL_26_DFFSR_70 gnd vdd FILL
XFILL_26_DFFSR_81 gnd vdd FILL
XFILL_26_DFFSR_92 gnd vdd FILL
XFILL_40_DFFSR_208 gnd vdd FILL
XFILL_8_AOI21X1_13 gnd vdd FILL
XFILL_40_DFFSR_219 gnd vdd FILL
XFILL_2_OAI21X1_9 gnd vdd FILL
XFILL_8_AOI21X1_24 gnd vdd FILL
XFILL_1_MUX2X1_1 gnd vdd FILL
XFILL_8_AOI21X1_35 gnd vdd FILL
XFILL_8_AOI21X1_46 gnd vdd FILL
XFILL_8_AOI21X1_57 gnd vdd FILL
XFILL_8_AOI21X1_68 gnd vdd FILL
XFILL_25_CLKBUF1_1 gnd vdd FILL
XFILL_18_OAI22X1_15 gnd vdd FILL
XFILL_18_OAI22X1_26 gnd vdd FILL
XFILL_66_DFFSR_80 gnd vdd FILL
XFILL_8_AOI21X1_79 gnd vdd FILL
XFILL_18_OAI22X1_37 gnd vdd FILL
XFILL_44_DFFSR_207 gnd vdd FILL
XFILL_66_DFFSR_91 gnd vdd FILL
XFILL_3_NOR2X1_11 gnd vdd FILL
XFILL_18_OAI22X1_48 gnd vdd FILL
XFILL_3_NOR2X1_22 gnd vdd FILL
XFILL_6_OAI21X1_8 gnd vdd FILL
XFILL_3_NOR2X1_33 gnd vdd FILL
XFILL_44_DFFSR_218 gnd vdd FILL
XFILL_3_NOR2X1_44 gnd vdd FILL
XFILL_44_DFFSR_229 gnd vdd FILL
XFILL_29_DFFSR_1 gnd vdd FILL
XFILL_3_NOR2X1_55 gnd vdd FILL
XFILL_2_CLKBUF1_16 gnd vdd FILL
XFILL_3_NOR2X1_66 gnd vdd FILL
XFILL_3_NOR2X1_77 gnd vdd FILL
XFILL_86_DFFSR_2 gnd vdd FILL
XFILL_3_NOR2X1_88 gnd vdd FILL
XFILL_2_CLKBUF1_27 gnd vdd FILL
XNAND3X1_90 NAND3X1_90/A NOR2X1_73/Y NOR3X1_25/Y gnd NOR2X1_74/A vdd NAND3X1
XFILL_2_CLKBUF1_38 gnd vdd FILL
XFILL_9_DFFSR_60 gnd vdd FILL
XFILL_3_NOR2X1_99 gnd vdd FILL
XFILL_7_NOR2X1_10 gnd vdd FILL
XFILL_48_DFFSR_206 gnd vdd FILL
XFILL_71_DFFSR_107 gnd vdd FILL
XFILL_9_DFFSR_71 gnd vdd FILL
XFILL_9_DFFSR_82 gnd vdd FILL
XFILL_48_DFFSR_217 gnd vdd FILL
XFILL_71_DFFSR_118 gnd vdd FILL
XFILL_7_NOR2X1_21 gnd vdd FILL
XFILL_9_DFFSR_93 gnd vdd FILL
XFILL_71_DFFSR_129 gnd vdd FILL
XFILL_7_NOR2X1_32 gnd vdd FILL
XFILL_7_NOR2X1_43 gnd vdd FILL
XFILL_48_DFFSR_228 gnd vdd FILL
XFILL_7_NOR2X1_54 gnd vdd FILL
XFILL_35_6_1 gnd vdd FILL
XFILL_48_DFFSR_239 gnd vdd FILL
XFILL_35_DFFSR_90 gnd vdd FILL
XFILL_11_OAI22X1_5 gnd vdd FILL
XFILL_7_NOR2X1_65 gnd vdd FILL
XFILL_34_1_0 gnd vdd FILL
XNOR2X1_90 NOR2X1_90/A NOR2X1_90/B gnd NOR2X1_90/Y vdd NOR2X1
XFILL_7_NOR2X1_76 gnd vdd FILL
XFILL_7_NOR2X1_87 gnd vdd FILL
XFILL_7_NOR2X1_98 gnd vdd FILL
XFILL_75_DFFSR_106 gnd vdd FILL
XFILL_0_NOR2X1_101 gnd vdd FILL
XFILL_11_OAI21X1_17 gnd vdd FILL
XFILL_75_DFFSR_117 gnd vdd FILL
XFILL_0_NOR2X1_112 gnd vdd FILL
XFILL_0_NOR2X1_123 gnd vdd FILL
XFILL_75_DFFSR_128 gnd vdd FILL
XFILL_0_NOR2X1_134 gnd vdd FILL
XFILL_11_OAI21X1_28 gnd vdd FILL
XFILL_75_DFFSR_139 gnd vdd FILL
XFILL_0_DFFSR_9 gnd vdd FILL
XFILL_0_NOR2X1_145 gnd vdd FILL
XFILL_15_OAI22X1_4 gnd vdd FILL
XFILL_11_OAI21X1_39 gnd vdd FILL
XFILL_0_NOR2X1_156 gnd vdd FILL
XFILL_13_DFFSR_7 gnd vdd FILL
XFILL_0_NOR2X1_167 gnd vdd FILL
XFILL_70_DFFSR_8 gnd vdd FILL
XFILL_0_NOR2X1_178 gnd vdd FILL
XFILL_79_DFFSR_105 gnd vdd FILL
XFILL_0_NOR2X1_189 gnd vdd FILL
XFILL_79_DFFSR_116 gnd vdd FILL
XFILL_79_DFFSR_127 gnd vdd FILL
XFILL_79_DFFSR_138 gnd vdd FILL
XFILL_79_DFFSR_149 gnd vdd FILL
XFILL_10_NAND2X1_60 gnd vdd FILL
XFILL_19_OAI22X1_3 gnd vdd FILL
XFILL_8_OAI22X1_10 gnd vdd FILL
XFILL_10_NAND2X1_71 gnd vdd FILL
XFILL_10_NAND2X1_82 gnd vdd FILL
XFILL_8_OAI22X1_21 gnd vdd FILL
XFILL_8_OAI22X1_32 gnd vdd FILL
XFILL_10_NAND2X1_93 gnd vdd FILL
XFILL_8_OAI22X1_43 gnd vdd FILL
XBUFX2_6 INVX2_3/A gnd addr[2] vdd BUFX2
XFILL_33_DFFSR_250 gnd vdd FILL
XFILL_33_DFFSR_261 gnd vdd FILL
XFILL_0_MUX2X1_107 gnd vdd FILL
XFILL_33_DFFSR_272 gnd vdd FILL
XFILL_0_MUX2X1_118 gnd vdd FILL
XFILL_0_MUX2X1_129 gnd vdd FILL
XFILL_5_NOR2X1_201 gnd vdd FILL
XFILL_60_DFFSR_150 gnd vdd FILL
XFILL_60_DFFSR_161 gnd vdd FILL
XFILL_37_DFFSR_260 gnd vdd FILL
XFILL_37_DFFSR_271 gnd vdd FILL
XFILL_60_DFFSR_172 gnd vdd FILL
XNAND2X1_1 NOR2X1_1/Y NOR2X1_13/Y gnd NOR2X1_57/A vdd NAND2X1
XFILL_60_DFFSR_183 gnd vdd FILL
XFILL_1_OAI21X1_12 gnd vdd FILL
XFILL_60_DFFSR_194 gnd vdd FILL
XFILL_7_NAND2X1_9 gnd vdd FILL
XFILL_1_OAI21X1_23 gnd vdd FILL
XFILL_3_MUX2X1_40 gnd vdd FILL
XFILL_1_OAI21X1_34 gnd vdd FILL
XFILL_11_DFFSR_207 gnd vdd FILL
XFILL_3_MUX2X1_51 gnd vdd FILL
XFILL_1_OAI21X1_45 gnd vdd FILL
XFILL_19_CLKBUF1_30 gnd vdd FILL
XFILL_11_DFFSR_218 gnd vdd FILL
XFILL_19_CLKBUF1_41 gnd vdd FILL
XFILL_3_MUX2X1_62 gnd vdd FILL
XFILL_11_DFFSR_229 gnd vdd FILL
XFILL_3_MUX2X1_73 gnd vdd FILL
XFILL_3_MUX2X1_84 gnd vdd FILL
XFILL_64_DFFSR_160 gnd vdd FILL
XFILL_3_MUX2X1_95 gnd vdd FILL
XFILL_64_DFFSR_171 gnd vdd FILL
XFILL_64_DFFSR_182 gnd vdd FILL
XFILL_64_DFFSR_193 gnd vdd FILL
XFILL_26_6_1 gnd vdd FILL
XFILL_15_DFFSR_206 gnd vdd FILL
XFILL_1_6_1 gnd vdd FILL
XFILL_14_AOI21X1_60 gnd vdd FILL
XFILL_14_AOI21X1_71 gnd vdd FILL
XFILL_12_NAND3X1_6 gnd vdd FILL
XFILL_7_MUX2X1_50 gnd vdd FILL
XFILL_15_DFFSR_217 gnd vdd FILL
XFILL_0_1_0 gnd vdd FILL
XFILL_7_MUX2X1_61 gnd vdd FILL
XFILL_25_1_0 gnd vdd FILL
XFILL_15_DFFSR_228 gnd vdd FILL
XFILL_15_DFFSR_239 gnd vdd FILL
XFILL_7_MUX2X1_72 gnd vdd FILL
XFILL_7_MUX2X1_83 gnd vdd FILL
XFILL_7_MUX2X1_94 gnd vdd FILL
XFILL_68_DFFSR_170 gnd vdd FILL
XNOR2X1_180 DFFSR_30/Q NOR2X1_181/B gnd NOR2X1_180/Y vdd NOR2X1
XNOR2X1_191 NOR2X1_68/A NOR2X1_7/B gnd NOR2X1_195/B vdd NOR2X1
XFILL_68_DFFSR_181 gnd vdd FILL
XFILL_68_DFFSR_192 gnd vdd FILL
XFILL_42_DFFSR_106 gnd vdd FILL
XFILL_19_DFFSR_205 gnd vdd FILL
XFILL_12_AND2X2_8 gnd vdd FILL
XFILL_19_DFFSR_216 gnd vdd FILL
XFILL_42_DFFSR_117 gnd vdd FILL
XFILL_42_DFFSR_128 gnd vdd FILL
XFILL_19_DFFSR_227 gnd vdd FILL
XFILL_42_DFFSR_139 gnd vdd FILL
XFILL_19_DFFSR_238 gnd vdd FILL
XFILL_19_DFFSR_249 gnd vdd FILL
XFILL_46_DFFSR_105 gnd vdd FILL
XAOI21X1_6 BUFX4_76/Y AOI21X1_7/B AOI21X1_6/C gnd DFFSR_141/D vdd AOI21X1
XFILL_46_DFFSR_116 gnd vdd FILL
XFILL_46_DFFSR_127 gnd vdd FILL
XFILL_46_DFFSR_138 gnd vdd FILL
XFILL_46_DFFSR_149 gnd vdd FILL
XMUX2X1_120 INVX1_162/Y BUFX4_76/Y NAND2X1_78/Y gnd DFFSR_137/D vdd MUX2X1
XMUX2X1_131 INVX1_175/Y MUX2X1_4/B NAND2X1_2/Y gnd DFFSR_121/D vdd MUX2X1
XMUX2X1_142 INVX1_186/Y BUFX4_72/Y NAND3X1_1/Y gnd DFFSR_115/D vdd MUX2X1
XMUX2X1_153 BUFX4_83/Y INVX1_197/Y NOR2X1_155/Y gnd DFFSR_89/D vdd MUX2X1
XFILL_17_MUX2X1_110 gnd vdd FILL
XMUX2X1_164 BUFX4_74/Y INVX1_209/Y NOR2X1_162/Y gnd DFFSR_78/D vdd MUX2X1
XFILL_17_MUX2X1_121 gnd vdd FILL
XMUX2X1_175 BUFX4_87/Y INVX1_220/Y NOR2X1_166/Y gnd DFFSR_63/D vdd MUX2X1
XFILL_17_MUX2X1_132 gnd vdd FILL
XMUX2X1_186 BUFX4_72/Y INVX1_5/Y NOR2X1_168/Y gnd DFFSR_56/D vdd MUX2X1
XFILL_23_MUX2X1_70 gnd vdd FILL
XFILL_17_MUX2X1_143 gnd vdd FILL
XFILL_9_7_1 gnd vdd FILL
XFILL_23_MUX2X1_81 gnd vdd FILL
XFILL_17_MUX2X1_154 gnd vdd FILL
XFILL_23_MUX2X1_92 gnd vdd FILL
XFILL_8_2_0 gnd vdd FILL
XFILL_17_MUX2X1_165 gnd vdd FILL
XFILL_17_MUX2X1_176 gnd vdd FILL
XFILL_17_MUX2X1_187 gnd vdd FILL
XINVX1_60 INVX1_60/A gnd INVX1_60/Y vdd INVX1
XFILL_30_DFFSR_1 gnd vdd FILL
XINVX1_71 INVX1_71/A gnd INVX1_71/Y vdd INVX1
XINVX1_82 INVX1_82/A gnd INVX1_82/Y vdd INVX1
XINVX1_93 INVX1_93/A gnd INVX1_93/Y vdd INVX1
XFILL_3_INVX1_15 gnd vdd FILL
XFILL_3_INVX1_26 gnd vdd FILL
XFILL_3_INVX1_37 gnd vdd FILL
XFILL_17_6_1 gnd vdd FILL
XFILL_31_DFFSR_160 gnd vdd FILL
XFILL_3_INVX1_48 gnd vdd FILL
XFILL_4_AND2X2_7 gnd vdd FILL
XFILL_3_INVX1_59 gnd vdd FILL
XFILL_16_1_0 gnd vdd FILL
XFILL_31_DFFSR_171 gnd vdd FILL
XFILL_31_DFFSR_182 gnd vdd FILL
XFILL_31_DFFSR_193 gnd vdd FILL
XFILL_49_DFFSR_18 gnd vdd FILL
XFILL_49_DFFSR_29 gnd vdd FILL
XFILL_35_DFFSR_170 gnd vdd FILL
XFILL_35_DFFSR_181 gnd vdd FILL
XFILL_35_DFFSR_192 gnd vdd FILL
XFILL_1_BUFX4_13 gnd vdd FILL
XFILL_52_DFFSR_5 gnd vdd FILL
XFILL_1_BUFX4_24 gnd vdd FILL
XFILL_1_BUFX4_35 gnd vdd FILL
XFILL_18_DFFSR_17 gnd vdd FILL
XFILL_1_BUFX4_46 gnd vdd FILL
XFILL_1_BUFX4_57 gnd vdd FILL
XFILL_7_MUX2X1_160 gnd vdd FILL
XFILL_1_BUFX4_68 gnd vdd FILL
XFILL_7_MUX2X1_171 gnd vdd FILL
XFILL_18_DFFSR_28 gnd vdd FILL
XFILL_18_DFFSR_39 gnd vdd FILL
XFILL_1_BUFX4_79 gnd vdd FILL
XFILL_39_DFFSR_180 gnd vdd FILL
XFILL_7_MUX2X1_182 gnd vdd FILL
XFILL_39_DFFSR_191 gnd vdd FILL
XFILL_7_MUX2X1_193 gnd vdd FILL
XFILL_13_DFFSR_105 gnd vdd FILL
XFILL_13_DFFSR_116 gnd vdd FILL
XFILL_13_DFFSR_127 gnd vdd FILL
XFILL_13_DFFSR_138 gnd vdd FILL
XFILL_58_DFFSR_16 gnd vdd FILL
XFILL_13_DFFSR_149 gnd vdd FILL
XFILL_58_DFFSR_27 gnd vdd FILL
XNOR2X1_4 NOR2X1_4/A NOR2X1_6/B gnd NOR2X1_4/Y vdd NOR2X1
XFILL_58_DFFSR_38 gnd vdd FILL
XFILL_58_DFFSR_49 gnd vdd FILL
XFILL_81_DFFSR_260 gnd vdd FILL
XFILL_17_DFFSR_104 gnd vdd FILL
XFILL_81_DFFSR_271 gnd vdd FILL
XFILL_17_DFFSR_115 gnd vdd FILL
XFILL_17_DFFSR_126 gnd vdd FILL
XFILL_17_DFFSR_137 gnd vdd FILL
XFILL_17_DFFSR_148 gnd vdd FILL
XFILL_17_DFFSR_8 gnd vdd FILL
XFILL_17_DFFSR_159 gnd vdd FILL
XFILL_74_DFFSR_9 gnd vdd FILL
XFILL_85_DFFSR_270 gnd vdd FILL
XFILL_27_DFFSR_15 gnd vdd FILL
XFILL_66_1 gnd vdd FILL
XFILL_27_DFFSR_26 gnd vdd FILL
XFILL_27_DFFSR_37 gnd vdd FILL
XFILL_66_0_0 gnd vdd FILL
XFILL_27_DFFSR_48 gnd vdd FILL
XFILL_27_DFFSR_59 gnd vdd FILL
XFILL_13_NOR3X1_16 gnd vdd FILL
XFILL_67_DFFSR_14 gnd vdd FILL
XFILL_13_NOR3X1_27 gnd vdd FILL
XFILL_67_DFFSR_25 gnd vdd FILL
XFILL_67_DFFSR_36 gnd vdd FILL
XFILL_13_NOR3X1_38 gnd vdd FILL
XFILL_13_NOR3X1_49 gnd vdd FILL
XFILL_63_DFFSR_205 gnd vdd FILL
XFILL_67_DFFSR_47 gnd vdd FILL
XFILL_67_DFFSR_58 gnd vdd FILL
XFILL_63_DFFSR_216 gnd vdd FILL
XFILL_63_DFFSR_227 gnd vdd FILL
XFILL_67_DFFSR_69 gnd vdd FILL
XFILL_63_DFFSR_238 gnd vdd FILL
XFILL_63_DFFSR_249 gnd vdd FILL
XFILL_17_NOR3X1_15 gnd vdd FILL
XFILL_17_NOR3X1_26 gnd vdd FILL
XFILL_50_4_1 gnd vdd FILL
XFILL_17_NOR3X1_37 gnd vdd FILL
XFILL_17_NOR3X1_48 gnd vdd FILL
XFILL_67_DFFSR_204 gnd vdd FILL
XFILL_67_DFFSR_215 gnd vdd FILL
XFILL_36_DFFSR_13 gnd vdd FILL
XFILL_36_DFFSR_24 gnd vdd FILL
XFILL_67_DFFSR_226 gnd vdd FILL
XFILL_36_DFFSR_35 gnd vdd FILL
XFILL_67_DFFSR_237 gnd vdd FILL
XFILL_36_DFFSR_46 gnd vdd FILL
XFILL_67_DFFSR_248 gnd vdd FILL
XFILL_36_DFFSR_57 gnd vdd FILL
XFILL_67_DFFSR_259 gnd vdd FILL
XFILL_36_DFFSR_68 gnd vdd FILL
XFILL_36_DFFSR_79 gnd vdd FILL
XAOI21X1_14 MUX2X1_1/A NOR2X1_153/B NOR2X1_150/Y gnd DFFSR_99/D vdd AOI21X1
XFILL_76_DFFSR_12 gnd vdd FILL
XAOI21X1_25 BUFX4_65/Y NOR2X1_181/B NOR2X1_179/Y gnd DFFSR_29/D vdd AOI21X1
XAOI21X1_36 BUFX4_65/Y NOR2X1_195/B NOR2X1_193/Y gnd DFFSR_16/D vdd AOI21X1
XAOI21X1_47 BUFX4_63/Y NOR2X1_6/B NOR2X1_4/Y gnd DFFSR_272/D vdd AOI21X1
XFILL_76_DFFSR_23 gnd vdd FILL
XFILL_76_DFFSR_34 gnd vdd FILL
XAOI21X1_58 BUFX4_97/Y NOR2X1_19/B NOR2X1_19/Y gnd DFFSR_257/D vdd AOI21X1
XFILL_3_NAND2X1_10 gnd vdd FILL
XFILL_76_DFFSR_45 gnd vdd FILL
XFILL_76_DFFSR_56 gnd vdd FILL
XAOI21X1_69 INVX1_126/Y INVX1_96/A OAI22X1_51/Y gnd NAND3X1_65/B vdd AOI21X1
XFILL_19_MUX2X1_2 gnd vdd FILL
XFILL_3_NAND2X1_21 gnd vdd FILL
XFILL_76_DFFSR_67 gnd vdd FILL
XFILL_3_NAND2X1_32 gnd vdd FILL
XFILL_76_DFFSR_78 gnd vdd FILL
XFILL_3_NAND2X1_43 gnd vdd FILL
XFILL_76_DFFSR_89 gnd vdd FILL
XFILL_3_NAND2X1_54 gnd vdd FILL
XFILL_3_NAND2X1_65 gnd vdd FILL
XOAI21X1_9 INVX1_34/Y OAI21X1_9/B OAI21X1_9/C gnd OAI21X1_9/Y vdd OAI21X1
XFILL_11_BUFX4_8 gnd vdd FILL
XFILL_3_NAND2X1_76 gnd vdd FILL
XFILL_3_NAND2X1_87 gnd vdd FILL
XFILL_45_DFFSR_11 gnd vdd FILL
XFILL_45_DFFSR_22 gnd vdd FILL
XFILL_45_DFFSR_33 gnd vdd FILL
XFILL_16_NOR3X1_8 gnd vdd FILL
XFILL_11_CLKBUF1_18 gnd vdd FILL
XFILL_45_DFFSR_44 gnd vdd FILL
XFILL_8_NOR2X1_19 gnd vdd FILL
XFILL_45_DFFSR_55 gnd vdd FILL
XFILL_11_CLKBUF1_29 gnd vdd FILL
XFILL_45_DFFSR_66 gnd vdd FILL
XFILL_45_DFFSR_77 gnd vdd FILL
XFILL_58_5_1 gnd vdd FILL
XFILL_45_DFFSR_88 gnd vdd FILL
XFILL_45_DFFSR_99 gnd vdd FILL
XFILL_85_DFFSR_10 gnd vdd FILL
XFILL_57_0_0 gnd vdd FILL
XFILL_85_DFFSR_21 gnd vdd FILL
XFILL_52_DFFSR_270 gnd vdd FILL
XFILL_85_DFFSR_32 gnd vdd FILL
XFILL_85_DFFSR_43 gnd vdd FILL
XFILL_14_DFFSR_10 gnd vdd FILL
XFILL_85_DFFSR_54 gnd vdd FILL
XFILL_29_CLKBUF1_20 gnd vdd FILL
XFILL_14_DFFSR_21 gnd vdd FILL
XFILL_85_DFFSR_65 gnd vdd FILL
XFILL_85_DFFSR_76 gnd vdd FILL
XFILL_29_CLKBUF1_31 gnd vdd FILL
XFILL_14_DFFSR_32 gnd vdd FILL
XFILL_85_DFFSR_87 gnd vdd FILL
XFILL_29_CLKBUF1_42 gnd vdd FILL
XFILL_14_DFFSR_43 gnd vdd FILL
XFILL_85_DFFSR_98 gnd vdd FILL
XFILL_14_DFFSR_54 gnd vdd FILL
XFILL_14_DFFSR_65 gnd vdd FILL
XFILL_14_DFFSR_76 gnd vdd FILL
XFILL_14_DFFSR_87 gnd vdd FILL
XFILL_30_DFFSR_205 gnd vdd FILL
XFILL_14_DFFSR_98 gnd vdd FILL
XFILL_7_AOI21X1_10 gnd vdd FILL
XFILL_54_DFFSR_20 gnd vdd FILL
XOAI22X1_11 INVX1_184/Y OAI22X1_50/B INVX1_180/Y OAI22X1_50/D gnd NOR2X1_64/B vdd
+ OAI22X1
XFILL_7_AOI21X1_21 gnd vdd FILL
XFILL_30_DFFSR_216 gnd vdd FILL
XFILL_54_DFFSR_31 gnd vdd FILL
XFILL_25_NOR3X1_6 gnd vdd FILL
XFILL_30_DFFSR_227 gnd vdd FILL
XFILL_54_DFFSR_42 gnd vdd FILL
XOAI22X1_22 INVX1_213/Y OAI22X1_48/B INVX1_217/Y OAI22X1_48/D gnd NOR2X1_82/A vdd
+ OAI22X1
XFILL_41_4_1 gnd vdd FILL
XFILL_7_AOI21X1_32 gnd vdd FILL
XFILL_30_DFFSR_238 gnd vdd FILL
XOAI22X1_33 INVX1_58/Y OAI22X1_33/B INVX1_62/Y OAI22X1_33/D gnd NOR2X1_96/B vdd OAI22X1
XFILL_7_AOI21X1_43 gnd vdd FILL
XOAI22X1_44 INVX1_112/Y OAI22X1_4/B MUX2X1_2/B OAI22X1_4/D gnd OAI22X1_44/Y vdd OAI22X1
XFILL_30_DFFSR_249 gnd vdd FILL
XFILL_54_DFFSR_53 gnd vdd FILL
XFILL_7_AOI21X1_54 gnd vdd FILL
XFILL_54_DFFSR_64 gnd vdd FILL
XFILL_54_DFFSR_75 gnd vdd FILL
XFILL_17_OAI22X1_12 gnd vdd FILL
XFILL_7_AOI21X1_65 gnd vdd FILL
XFILL_83_DFFSR_180 gnd vdd FILL
XFILL_54_DFFSR_86 gnd vdd FILL
XFILL_17_OAI22X1_23 gnd vdd FILL
XFILL_17_OAI22X1_34 gnd vdd FILL
XFILL_7_AOI21X1_76 gnd vdd FILL
XFILL_83_DFFSR_191 gnd vdd FILL
XFILL_54_DFFSR_97 gnd vdd FILL
XFILL_34_DFFSR_204 gnd vdd FILL
XFILL_17_OAI22X1_45 gnd vdd FILL
XFILL_34_DFFSR_215 gnd vdd FILL
XFILL_34_DFFSR_226 gnd vdd FILL
XFILL_34_DFFSR_237 gnd vdd FILL
XFILL_34_DFFSR_2 gnd vdd FILL
XFILL_3_DFFSR_250 gnd vdd FILL
XFILL_34_DFFSR_248 gnd vdd FILL
XFILL_3_DFFSR_261 gnd vdd FILL
XFILL_3_DFFSR_272 gnd vdd FILL
XFILL_1_CLKBUF1_13 gnd vdd FILL
XFILL_34_DFFSR_259 gnd vdd FILL
XFILL_1_CLKBUF1_24 gnd vdd FILL
XFILL_23_DFFSR_30 gnd vdd FILL
XFILL_23_DFFSR_41 gnd vdd FILL
XFILL_0_MUX2X1_17 gnd vdd FILL
XFILL_87_DFFSR_190 gnd vdd FILL
XFILL_1_CLKBUF1_35 gnd vdd FILL
XFILL_23_DFFSR_52 gnd vdd FILL
XFILL_0_MUX2X1_28 gnd vdd FILL
XFILL_61_DFFSR_104 gnd vdd FILL
XFILL_0_MUX2X1_39 gnd vdd FILL
XFILL_38_DFFSR_203 gnd vdd FILL
XFILL_23_DFFSR_63 gnd vdd FILL
XFILL_61_DFFSR_115 gnd vdd FILL
XFILL_38_DFFSR_214 gnd vdd FILL
XFILL_23_DFFSR_74 gnd vdd FILL
XFILL_61_DFFSR_126 gnd vdd FILL
XFILL_38_DFFSR_225 gnd vdd FILL
XFILL_61_DFFSR_137 gnd vdd FILL
XFILL_23_DFFSR_85 gnd vdd FILL
XFILL_61_DFFSR_148 gnd vdd FILL
XFILL_23_DFFSR_96 gnd vdd FILL
XFILL_38_DFFSR_236 gnd vdd FILL
XFILL_38_DFFSR_247 gnd vdd FILL
XFILL_7_DFFSR_260 gnd vdd FILL
XFILL_8_NOR3X1_7 gnd vdd FILL
XFILL_7_DFFSR_271 gnd vdd FILL
XFILL_38_DFFSR_258 gnd vdd FILL
XFILL_61_DFFSR_159 gnd vdd FILL
XFILL_38_DFFSR_269 gnd vdd FILL
XFILL_63_DFFSR_40 gnd vdd FILL
XFILL_4_MUX2X1_16 gnd vdd FILL
XFILL_63_DFFSR_51 gnd vdd FILL
XFILL_65_DFFSR_103 gnd vdd FILL
XFILL_4_MUX2X1_27 gnd vdd FILL
XFILL_63_DFFSR_62 gnd vdd FILL
XFILL_4_MUX2X1_38 gnd vdd FILL
XFILL_10_OAI21X1_14 gnd vdd FILL
XFILL_65_DFFSR_114 gnd vdd FILL
XFILL_4_MUX2X1_49 gnd vdd FILL
XFILL_10_OAI21X1_25 gnd vdd FILL
XFILL_63_DFFSR_73 gnd vdd FILL
XFILL_65_DFFSR_125 gnd vdd FILL
XFILL_65_DFFSR_136 gnd vdd FILL
XFILL_63_DFFSR_84 gnd vdd FILL
XFILL_63_DFFSR_95 gnd vdd FILL
XFILL_10_OAI21X1_36 gnd vdd FILL
XFILL_65_DFFSR_147 gnd vdd FILL
XFILL_10_OAI21X1_47 gnd vdd FILL
XFILL_65_DFFSR_158 gnd vdd FILL
XFILL_65_DFFSR_169 gnd vdd FILL
XFILL_6_DFFSR_20 gnd vdd FILL
XFILL_8_MUX2X1_15 gnd vdd FILL
XFILL_69_DFFSR_102 gnd vdd FILL
XFILL_6_DFFSR_31 gnd vdd FILL
XFILL_8_MUX2X1_26 gnd vdd FILL
XFILL_49_5_1 gnd vdd FILL
XFILL_8_MUX2X1_37 gnd vdd FILL
XFILL_6_DFFSR_42 gnd vdd FILL
XFILL_56_DFFSR_6 gnd vdd FILL
XFILL_8_MUX2X1_48 gnd vdd FILL
XFILL_6_DFFSR_53 gnd vdd FILL
XFILL_69_DFFSR_113 gnd vdd FILL
XFILL_69_DFFSR_124 gnd vdd FILL
XFILL_8_MUX2X1_59 gnd vdd FILL
XFILL_48_0_0 gnd vdd FILL
XFILL_69_DFFSR_135 gnd vdd FILL
XFILL_6_DFFSR_64 gnd vdd FILL
XFILL_69_DFFSR_146 gnd vdd FILL
XFILL_12_OAI21X1_3 gnd vdd FILL
XFILL_6_DFFSR_75 gnd vdd FILL
XFILL_32_DFFSR_50 gnd vdd FILL
XFILL_69_DFFSR_157 gnd vdd FILL
XFILL_6_DFFSR_86 gnd vdd FILL
XFILL_32_DFFSR_61 gnd vdd FILL
XFILL_32_DFFSR_72 gnd vdd FILL
XFILL_6_DFFSR_97 gnd vdd FILL
XFILL_69_DFFSR_168 gnd vdd FILL
XFILL_32_DFFSR_83 gnd vdd FILL
XFILL_69_DFFSR_179 gnd vdd FILL
XFILL_7_OAI22X1_40 gnd vdd FILL
XFILL_7_OAI22X1_51 gnd vdd FILL
XFILL_32_DFFSR_94 gnd vdd FILL
XFILL_0_INVX1_210 gnd vdd FILL
XFILL_0_INVX1_221 gnd vdd FILL
XFILL_38_5 gnd vdd FILL
XFILL_72_DFFSR_60 gnd vdd FILL
XFILL_72_DFFSR_71 gnd vdd FILL
XFILL_72_DFFSR_82 gnd vdd FILL
XFILL_72_DFFSR_93 gnd vdd FILL
XFILL_20_MUX2X1_14 gnd vdd FILL
XFILL_32_4_1 gnd vdd FILL
XFILL_4_INVX1_220 gnd vdd FILL
XFILL_20_MUX2X1_25 gnd vdd FILL
XFILL_20_MUX2X1_36 gnd vdd FILL
XFILL_20_MUX2X1_47 gnd vdd FILL
XFILL_20_MUX2X1_58 gnd vdd FILL
XFILL_20_MUX2X1_69 gnd vdd FILL
XFILL_12_NOR3X1_1 gnd vdd FILL
XFILL_50_DFFSR_180 gnd vdd FILL
XFILL_0_OAI21X1_20 gnd vdd FILL
XFILL_50_DFFSR_191 gnd vdd FILL
XFILL_0_OAI21X1_31 gnd vdd FILL
XFILL_41_DFFSR_70 gnd vdd FILL
XFILL_41_DFFSR_81 gnd vdd FILL
XFILL_0_OAI21X1_42 gnd vdd FILL
XFILL_41_DFFSR_92 gnd vdd FILL
XFILL_54_DFFSR_190 gnd vdd FILL
XFILL_81_DFFSR_80 gnd vdd FILL
XFILL_81_DFFSR_91 gnd vdd FILL
XFILL_10_DFFSR_80 gnd vdd FILL
XFILL_10_DFFSR_91 gnd vdd FILL
XFILL_32_DFFSR_103 gnd vdd FILL
XFILL_32_DFFSR_114 gnd vdd FILL
XFILL_32_DFFSR_125 gnd vdd FILL
XFILL_32_DFFSR_136 gnd vdd FILL
XFILL_32_DFFSR_147 gnd vdd FILL
XFILL_1_DFFSR_160 gnd vdd FILL
XFILL_21_10 gnd vdd FILL
XFILL_32_DFFSR_158 gnd vdd FILL
XFILL_1_DFFSR_171 gnd vdd FILL
XFILL_50_DFFSR_90 gnd vdd FILL
XFILL_32_DFFSR_169 gnd vdd FILL
XFILL_1_DFFSR_182 gnd vdd FILL
XFILL_39_0_0 gnd vdd FILL
XFILL_1_DFFSR_193 gnd vdd FILL
XFILL_36_DFFSR_102 gnd vdd FILL
XFILL_36_DFFSR_113 gnd vdd FILL
XFILL_36_DFFSR_124 gnd vdd FILL
XFILL_2_NAND3X1_18 gnd vdd FILL
XFILL_36_DFFSR_135 gnd vdd FILL
XFILL_2_NAND3X1_29 gnd vdd FILL
XFILL_36_DFFSR_146 gnd vdd FILL
XFILL_36_DFFSR_157 gnd vdd FILL
XFILL_5_DFFSR_170 gnd vdd FILL
XFILL_36_DFFSR_168 gnd vdd FILL
XFILL_5_DFFSR_181 gnd vdd FILL
XFILL_36_DFFSR_179 gnd vdd FILL
XFILL_5_DFFSR_192 gnd vdd FILL
XFILL_15_BUFX4_9 gnd vdd FILL
XFILL_16_MUX2X1_140 gnd vdd FILL
XFILL_23_4_1 gnd vdd FILL
XFILL_9_DFFSR_180 gnd vdd FILL
XFILL_16_MUX2X1_151 gnd vdd FILL
XFILL_16_MUX2X1_162 gnd vdd FILL
XFILL_9_DFFSR_191 gnd vdd FILL
XFILL_16_MUX2X1_173 gnd vdd FILL
XFILL_16_MUX2X1_184 gnd vdd FILL
XFILL_82_DFFSR_203 gnd vdd FILL
XFILL_82_DFFSR_214 gnd vdd FILL
XFILL_82_DFFSR_225 gnd vdd FILL
XFILL_82_DFFSR_236 gnd vdd FILL
XFILL_3_DFFSR_1 gnd vdd FILL
XFILL_82_DFFSR_247 gnd vdd FILL
XFILL_82_DFFSR_258 gnd vdd FILL
XFILL_82_DFFSR_269 gnd vdd FILL
XFILL_86_DFFSR_202 gnd vdd FILL
XFILL_86_DFFSR_213 gnd vdd FILL
XFILL_2_DFFSR_90 gnd vdd FILL
XFILL_86_DFFSR_224 gnd vdd FILL
XFILL_13_AOI21X1_9 gnd vdd FILL
XFILL_86_DFFSR_235 gnd vdd FILL
XFILL_86_DFFSR_246 gnd vdd FILL
XFILL_86_DFFSR_257 gnd vdd FILL
XFILL_86_DFFSR_268 gnd vdd FILL
XFILL_21_DFFSR_190 gnd vdd FILL
XFILL_11_BUFX2_5 gnd vdd FILL
XFILL_2_INVX1_130 gnd vdd FILL
XFILL_2_INVX1_141 gnd vdd FILL
XFILL_2_INVX1_152 gnd vdd FILL
XFILL_2_INVX1_163 gnd vdd FILL
XFILL_2_INVX1_174 gnd vdd FILL
XFILL_2_INVX1_185 gnd vdd FILL
XFILL_2_INVX1_196 gnd vdd FILL
XFILL_21_CLKBUF1_19 gnd vdd FILL
XFILL_6_5_1 gnd vdd FILL
XFILL_6_INVX1_140 gnd vdd FILL
XFILL_6_INVX1_151 gnd vdd FILL
XFILL_38_DFFSR_3 gnd vdd FILL
XFILL_6_INVX1_162 gnd vdd FILL
XFILL_5_0_0 gnd vdd FILL
XFILL_0_INVX1_19 gnd vdd FILL
XFILL_6_INVX1_173 gnd vdd FILL
XFILL_6_INVX1_184 gnd vdd FILL
XFILL_6_INVX1_195 gnd vdd FILL
XFILL_6_MUX2X1_190 gnd vdd FILL
XFILL_0_OAI22X1_3 gnd vdd FILL
XFILL_14_4_1 gnd vdd FILL
XFILL_2_NOR2X1_108 gnd vdd FILL
XFILL_2_NOR2X1_119 gnd vdd FILL
XFILL_4_OAI22X1_2 gnd vdd FILL
XFILL_22_DFFSR_9 gnd vdd FILL
XFILL_8_OAI22X1_1 gnd vdd FILL
XFILL_53_DFFSR_202 gnd vdd FILL
XFILL_53_DFFSR_213 gnd vdd FILL
XFILL_53_DFFSR_224 gnd vdd FILL
XFILL_53_DFFSR_235 gnd vdd FILL
XFILL_53_DFFSR_246 gnd vdd FILL
XFILL_53_DFFSR_257 gnd vdd FILL
XFILL_53_DFFSR_268 gnd vdd FILL
XFILL_9_NAND3X1_60 gnd vdd FILL
XFILL_9_NAND3X1_71 gnd vdd FILL
XFILL_9_NAND3X1_82 gnd vdd FILL
XFILL_57_DFFSR_201 gnd vdd FILL
XFILL_9_NAND3X1_93 gnd vdd FILL
XFILL_80_DFFSR_102 gnd vdd FILL
XFILL_24_DFFSR_19 gnd vdd FILL
XFILL_15_BUFX4_40 gnd vdd FILL
XFILL_57_DFFSR_212 gnd vdd FILL
XFILL_80_DFFSR_113 gnd vdd FILL
XFILL_80_DFFSR_124 gnd vdd FILL
XFILL_15_BUFX4_51 gnd vdd FILL
XFILL_57_DFFSR_223 gnd vdd FILL
XFILL_1_3 gnd vdd FILL
XFILL_80_DFFSR_135 gnd vdd FILL
XFILL_15_BUFX4_62 gnd vdd FILL
XFILL_80_DFFSR_146 gnd vdd FILL
XFILL_57_DFFSR_234 gnd vdd FILL
XFILL_15_BUFX4_73 gnd vdd FILL
XFILL_57_DFFSR_245 gnd vdd FILL
XFILL_80_DFFSR_157 gnd vdd FILL
XFILL_15_BUFX4_84 gnd vdd FILL
XFILL_57_DFFSR_256 gnd vdd FILL
XFILL_15_BUFX4_95 gnd vdd FILL
XFILL_57_DFFSR_267 gnd vdd FILL
XFILL_80_DFFSR_168 gnd vdd FILL
XFILL_80_DFFSR_179 gnd vdd FILL
XFILL_12_CLKBUF1_8 gnd vdd FILL
XFILL_12_AOI22X1_10 gnd vdd FILL
XFILL_0_DFFSR_205 gnd vdd FILL
XFILL_84_DFFSR_101 gnd vdd FILL
XFILL_3_OAI21X1_19 gnd vdd FILL
XFILL_0_DFFSR_216 gnd vdd FILL
XFILL_64_DFFSR_18 gnd vdd FILL
XFILL_84_DFFSR_112 gnd vdd FILL
XFILL_50_4 gnd vdd FILL
XFILL_0_DFFSR_227 gnd vdd FILL
XFILL_64_DFFSR_29 gnd vdd FILL
XFILL_84_DFFSR_123 gnd vdd FILL
XFILL_84_DFFSR_134 gnd vdd FILL
XFILL_0_DFFSR_238 gnd vdd FILL
XFILL_84_DFFSR_145 gnd vdd FILL
XFILL_0_DFFSR_249 gnd vdd FILL
XFILL_64_3_1 gnd vdd FILL
XFILL_84_DFFSR_156 gnd vdd FILL
XFILL_43_3 gnd vdd FILL
XFILL_84_DFFSR_167 gnd vdd FILL
XFILL_16_CLKBUF1_7 gnd vdd FILL
XFILL_84_DFFSR_178 gnd vdd FILL
XFILL_84_DFFSR_189 gnd vdd FILL
XFILL_2_NAND2X1_40 gnd vdd FILL
XFILL_4_DFFSR_204 gnd vdd FILL
XFILL_4_DFFSR_215 gnd vdd FILL
XFILL_2_NAND2X1_51 gnd vdd FILL
XFILL_1_NAND3X1_4 gnd vdd FILL
XFILL_2_NAND2X1_62 gnd vdd FILL
XFILL_2_NAND2X1_73 gnd vdd FILL
XFILL_4_DFFSR_226 gnd vdd FILL
XFILL_4_DFFSR_237 gnd vdd FILL
XFILL_4_DFFSR_248 gnd vdd FILL
XFILL_2_NAND2X1_84 gnd vdd FILL
XFILL_12_BUFX4_102 gnd vdd FILL
XFILL_2_NAND2X1_95 gnd vdd FILL
XFILL_4_DFFSR_259 gnd vdd FILL
XFILL_33_DFFSR_17 gnd vdd FILL
XFILL_33_DFFSR_28 gnd vdd FILL
XFILL_33_DFFSR_39 gnd vdd FILL
XFILL_8_DFFSR_203 gnd vdd FILL
XFILL_5_NAND3X1_3 gnd vdd FILL
XFILL_10_CLKBUF1_15 gnd vdd FILL
XFILL_8_DFFSR_214 gnd vdd FILL
XFILL_10_CLKBUF1_26 gnd vdd FILL
XFILL_8_DFFSR_225 gnd vdd FILL
XFILL_10_CLKBUF1_37 gnd vdd FILL
XFILL_8_DFFSR_236 gnd vdd FILL
XFILL_8_DFFSR_247 gnd vdd FILL
XFILL_73_DFFSR_16 gnd vdd FILL
XFILL_8_DFFSR_258 gnd vdd FILL
XFILL_8_DFFSR_269 gnd vdd FILL
XFILL_73_DFFSR_27 gnd vdd FILL
XFILL_73_DFFSR_38 gnd vdd FILL
XFILL_73_DFFSR_49 gnd vdd FILL
XFILL_9_NAND3X1_2 gnd vdd FILL
XFILL_16_MUX2X1_6 gnd vdd FILL
XFILL_16_10 gnd vdd FILL
XFILL_7_BUFX4_50 gnd vdd FILL
XFILL_7_BUFX4_61 gnd vdd FILL
XFILL_42_DFFSR_15 gnd vdd FILL
XFILL_20_DFFSR_202 gnd vdd FILL
XFILL_42_DFFSR_26 gnd vdd FILL
XFILL_7_BUFX4_72 gnd vdd FILL
XFILL_7_BUFX4_83 gnd vdd FILL
XFILL_20_DFFSR_213 gnd vdd FILL
XFILL_19_MUX2X1_106 gnd vdd FILL
XFILL_42_DFFSR_37 gnd vdd FILL
XFILL_10_NOR2X1_15 gnd vdd FILL
XFILL_7_BUFX4_94 gnd vdd FILL
XFILL_19_MUX2X1_117 gnd vdd FILL
XFILL_10_NOR2X1_26 gnd vdd FILL
XFILL_42_DFFSR_48 gnd vdd FILL
XFILL_1_AOI22X1_9 gnd vdd FILL
XFILL_20_DFFSR_224 gnd vdd FILL
XFILL_20_DFFSR_235 gnd vdd FILL
XFILL_10_NOR2X1_37 gnd vdd FILL
XFILL_19_MUX2X1_128 gnd vdd FILL
XFILL_42_DFFSR_59 gnd vdd FILL
XFILL_6_AOI21X1_40 gnd vdd FILL
XFILL_19_MUX2X1_139 gnd vdd FILL
XFILL_20_DFFSR_246 gnd vdd FILL
XFILL_10_NOR2X1_48 gnd vdd FILL
XFILL_6_AOI21X1_51 gnd vdd FILL
XFILL_20_DFFSR_257 gnd vdd FILL
XFILL_20_DFFSR_268 gnd vdd FILL
XFILL_10_NOR2X1_59 gnd vdd FILL
XFILL_6_AOI21X1_62 gnd vdd FILL
XFILL_6_AOI21X1_73 gnd vdd FILL
XFILL_16_OAI22X1_20 gnd vdd FILL
XFILL_1_INVX1_208 gnd vdd FILL
XFILL_16_OAI22X1_31 gnd vdd FILL
XFILL_82_DFFSR_14 gnd vdd FILL
XFILL_24_DFFSR_201 gnd vdd FILL
XFILL_16_OAI22X1_42 gnd vdd FILL
XFILL_82_DFFSR_25 gnd vdd FILL
XFILL_82_DFFSR_36 gnd vdd FILL
XFILL_24_DFFSR_212 gnd vdd FILL
XFILL_1_INVX1_219 gnd vdd FILL
XFILL_24_DFFSR_223 gnd vdd FILL
XFILL_5_AOI22X1_8 gnd vdd FILL
XFILL_82_DFFSR_47 gnd vdd FILL
XFILL_24_DFFSR_234 gnd vdd FILL
XFILL_82_DFFSR_58 gnd vdd FILL
XFILL_11_DFFSR_14 gnd vdd FILL
XFILL_7_DFFSR_2 gnd vdd FILL
XFILL_82_DFFSR_69 gnd vdd FILL
XFILL_11_DFFSR_25 gnd vdd FILL
XFILL_24_DFFSR_245 gnd vdd FILL
XFILL_9_NOR2X1_150 gnd vdd FILL
XFILL_11_DFFSR_36 gnd vdd FILL
XFILL_0_CLKBUF1_10 gnd vdd FILL
XFILL_24_DFFSR_256 gnd vdd FILL
XFILL_0_CLKBUF1_21 gnd vdd FILL
XFILL_9_NOR2X1_161 gnd vdd FILL
XFILL_24_DFFSR_267 gnd vdd FILL
XFILL_0_CLKBUF1_32 gnd vdd FILL
XFILL_11_DFFSR_47 gnd vdd FILL
XFILL_5_INVX1_207 gnd vdd FILL
XFILL_51_DFFSR_101 gnd vdd FILL
XFILL_11_DFFSR_58 gnd vdd FILL
XFILL_77_DFFSR_1 gnd vdd FILL
XFILL_9_NOR2X1_172 gnd vdd FILL
XFILL_28_DFFSR_200 gnd vdd FILL
XFILL_9_NOR2X1_7 gnd vdd FILL
XFILL_9_NOR2X1_183 gnd vdd FILL
XFILL_11_DFFSR_69 gnd vdd FILL
XFILL_5_INVX1_218 gnd vdd FILL
XFILL_28_DFFSR_211 gnd vdd FILL
XFILL_55_3_1 gnd vdd FILL
XFILL_9_NOR2X1_194 gnd vdd FILL
XFILL_51_DFFSR_112 gnd vdd FILL
XFILL_28_DFFSR_222 gnd vdd FILL
XFILL_51_DFFSR_123 gnd vdd FILL
XFILL_51_DFFSR_134 gnd vdd FILL
XFILL_28_DFFSR_233 gnd vdd FILL
XFILL_9_AOI22X1_7 gnd vdd FILL
XFILL_51_DFFSR_13 gnd vdd FILL
XFILL_51_DFFSR_145 gnd vdd FILL
XFILL_51_DFFSR_24 gnd vdd FILL
XFILL_28_DFFSR_244 gnd vdd FILL
XFILL_51_DFFSR_156 gnd vdd FILL
XFILL_51_DFFSR_35 gnd vdd FILL
XFILL_28_DFFSR_255 gnd vdd FILL
XFILL_2_BUFX2_8 gnd vdd FILL
XFILL_51_DFFSR_46 gnd vdd FILL
XFILL_51_DFFSR_167 gnd vdd FILL
XFILL_28_DFFSR_266 gnd vdd FILL
XFILL_51_DFFSR_178 gnd vdd FILL
XFILL_51_DFFSR_57 gnd vdd FILL
XFILL_55_DFFSR_100 gnd vdd FILL
XFILL_51_DFFSR_189 gnd vdd FILL
XFILL_51_DFFSR_68 gnd vdd FILL
XFILL_55_DFFSR_111 gnd vdd FILL
XFILL_51_DFFSR_79 gnd vdd FILL
XFILL_55_DFFSR_122 gnd vdd FILL
XFILL_55_DFFSR_133 gnd vdd FILL
XFILL_55_DFFSR_144 gnd vdd FILL
XFILL_55_DFFSR_155 gnd vdd FILL
XFILL_8_MUX2X1_5 gnd vdd FILL
XFILL_55_DFFSR_166 gnd vdd FILL
XFILL_55_DFFSR_177 gnd vdd FILL
XFILL_20_DFFSR_12 gnd vdd FILL
XFILL_55_DFFSR_188 gnd vdd FILL
XFILL_9_MUX2X1_101 gnd vdd FILL
XFILL_9_MUX2X1_112 gnd vdd FILL
XFILL_59_DFFSR_110 gnd vdd FILL
XFILL_55_DFFSR_199 gnd vdd FILL
XFILL_20_DFFSR_23 gnd vdd FILL
XFILL_61_DFFSR_7 gnd vdd FILL
XFILL_9_MUX2X1_123 gnd vdd FILL
XFILL_20_DFFSR_34 gnd vdd FILL
XFILL_59_DFFSR_121 gnd vdd FILL
XFILL_20_DFFSR_45 gnd vdd FILL
XFILL_9_MUX2X1_134 gnd vdd FILL
XFILL_20_DFFSR_56 gnd vdd FILL
XFILL_59_DFFSR_132 gnd vdd FILL
XFILL_9_MUX2X1_145 gnd vdd FILL
XFILL_59_DFFSR_143 gnd vdd FILL
XFILL_59_DFFSR_154 gnd vdd FILL
XFILL_9_MUX2X1_156 gnd vdd FILL
XFILL_20_DFFSR_67 gnd vdd FILL
XFILL_20_DFFSR_78 gnd vdd FILL
XFILL_59_DFFSR_165 gnd vdd FILL
XFILL_9_MUX2X1_167 gnd vdd FILL
XFILL_20_DFFSR_89 gnd vdd FILL
XFILL_9_MUX2X1_178 gnd vdd FILL
XFILL_60_DFFSR_11 gnd vdd FILL
XFILL_2_DFFSR_103 gnd vdd FILL
XFILL_59_DFFSR_176 gnd vdd FILL
XFILL_9_MUX2X1_189 gnd vdd FILL
XFILL_59_DFFSR_187 gnd vdd FILL
XFILL_59_DFFSR_198 gnd vdd FILL
XFILL_60_DFFSR_22 gnd vdd FILL
XFILL_2_DFFSR_114 gnd vdd FILL
XFILL_60_DFFSR_33 gnd vdd FILL
XFILL_2_DFFSR_125 gnd vdd FILL
XFILL_2_DFFSR_136 gnd vdd FILL
XFILL_31_NOR3X1_8 gnd vdd FILL
XFILL_60_DFFSR_44 gnd vdd FILL
XFILL_60_DFFSR_55 gnd vdd FILL
XFILL_2_DFFSR_147 gnd vdd FILL
XFILL_60_DFFSR_66 gnd vdd FILL
XFILL_2_DFFSR_158 gnd vdd FILL
XDFFSR_80 DFFSR_80/Q DFFSR_84/CLK DFFSR_84/R vdd DFFSR_80/D gnd vdd DFFSR
XFILL_60_DFFSR_77 gnd vdd FILL
XFILL_2_DFFSR_169 gnd vdd FILL
XDFFSR_91 DFFSR_91/Q CLKBUF1_1/Y DFFSR_91/R vdd DFFSR_91/D gnd vdd DFFSR
XFILL_60_DFFSR_88 gnd vdd FILL
XFILL_6_DFFSR_102 gnd vdd FILL
XFILL_60_DFFSR_99 gnd vdd FILL
XFILL_10_MUX2X1_11 gnd vdd FILL
XFILL_6_DFFSR_113 gnd vdd FILL
XFILL_6_DFFSR_124 gnd vdd FILL
XFILL_3_DFFSR_13 gnd vdd FILL
XFILL_10_MUX2X1_22 gnd vdd FILL
XFILL_3_DFFSR_24 gnd vdd FILL
XFILL_6_DFFSR_135 gnd vdd FILL
XFILL_10_MUX2X1_33 gnd vdd FILL
XFILL_6_DFFSR_146 gnd vdd FILL
XFILL_3_DFFSR_35 gnd vdd FILL
XFILL_1_BUFX4_2 gnd vdd FILL
XFILL_10_MUX2X1_44 gnd vdd FILL
XFILL_6_DFFSR_157 gnd vdd FILL
XFILL_3_DFFSR_46 gnd vdd FILL
XFILL_10_MUX2X1_55 gnd vdd FILL
XFILL_3_DFFSR_57 gnd vdd FILL
XFILL_10_MUX2X1_66 gnd vdd FILL
XFILL_6_DFFSR_168 gnd vdd FILL
XFILL_10_MUX2X1_77 gnd vdd FILL
XFILL_6_DFFSR_179 gnd vdd FILL
XFILL_3_DFFSR_68 gnd vdd FILL
XFILL_10_MUX2X1_88 gnd vdd FILL
XFILL_3_DFFSR_79 gnd vdd FILL
XFILL_10_MUX2X1_99 gnd vdd FILL
XFILL_14_MUX2X1_10 gnd vdd FILL
XFILL_14_MUX2X1_21 gnd vdd FILL
XFILL_14_MUX2X1_32 gnd vdd FILL
XFILL_14_MUX2X1_43 gnd vdd FILL
XFILL_14_MUX2X1_54 gnd vdd FILL
XFILL_14_MUX2X1_65 gnd vdd FILL
XFILL_2_NOR3X1_14 gnd vdd FILL
XFILL_14_MUX2X1_76 gnd vdd FILL
XFILL_46_3_1 gnd vdd FILL
XFILL_14_MUX2X1_87 gnd vdd FILL
XFILL_2_NOR3X1_25 gnd vdd FILL
XFILL_14_MUX2X1_98 gnd vdd FILL
XFILL_2_NOR3X1_36 gnd vdd FILL
XFILL_18_MUX2X1_20 gnd vdd FILL
XFILL_2_NOR3X1_47 gnd vdd FILL
XFILL_18_MUX2X1_31 gnd vdd FILL
XFILL_18_MUX2X1_42 gnd vdd FILL
XFILL_18_MUX2X1_53 gnd vdd FILL
XFILL_18_MUX2X1_64 gnd vdd FILL
XFILL_0_INVX1_6 gnd vdd FILL
XFILL_6_NOR3X1_13 gnd vdd FILL
XFILL_18_MUX2X1_75 gnd vdd FILL
XFILL_18_MUX2X1_86 gnd vdd FILL
XFILL_6_NOR3X1_24 gnd vdd FILL
XFILL_18_MUX2X1_97 gnd vdd FILL
XFILL_6_NOR3X1_35 gnd vdd FILL
XFILL_22_8 gnd vdd FILL
XFILL_22_DFFSR_100 gnd vdd FILL
XFILL_6_NOR3X1_46 gnd vdd FILL
XFILL_22_DFFSR_111 gnd vdd FILL
XFILL_22_DFFSR_122 gnd vdd FILL
XFILL_22_DFFSR_133 gnd vdd FILL
XFILL_30_7_2 gnd vdd FILL
XFILL_22_DFFSR_144 gnd vdd FILL
XFILL_22_DFFSR_155 gnd vdd FILL
XFILL_22_DFFSR_166 gnd vdd FILL
XFILL_22_DFFSR_177 gnd vdd FILL
XFILL_3_INVX1_106 gnd vdd FILL
XFILL_22_DFFSR_188 gnd vdd FILL
XFILL_3_INVX1_117 gnd vdd FILL
XFILL_26_DFFSR_110 gnd vdd FILL
XFILL_22_DFFSR_199 gnd vdd FILL
XFILL_3_INVX1_128 gnd vdd FILL
XFILL_1_NAND3X1_15 gnd vdd FILL
XFILL_3_INVX1_139 gnd vdd FILL
XFILL_26_DFFSR_121 gnd vdd FILL
XFILL_26_DFFSR_132 gnd vdd FILL
XFILL_1_NAND3X1_26 gnd vdd FILL
XFILL_26_DFFSR_143 gnd vdd FILL
XFILL_1_NAND3X1_37 gnd vdd FILL
XFILL_26_DFFSR_154 gnd vdd FILL
XFILL_1_NAND3X1_48 gnd vdd FILL
XFILL_26_DFFSR_165 gnd vdd FILL
XFILL_1_NAND3X1_59 gnd vdd FILL
XFILL_5_NAND2X1_17 gnd vdd FILL
XFILL_7_INVX1_105 gnd vdd FILL
XFILL_5_NAND2X1_28 gnd vdd FILL
XFILL_26_DFFSR_176 gnd vdd FILL
XFILL_26_DFFSR_187 gnd vdd FILL
XFILL_26_DFFSR_198 gnd vdd FILL
XFILL_7_INVX1_116 gnd vdd FILL
XINVX1_130 INVX1_130/A gnd INVX1_130/Y vdd INVX1
XFILL_5_NAND2X1_39 gnd vdd FILL
XFILL_7_INVX1_127 gnd vdd FILL
XINVX1_141 NOR2X1_24/A gnd INVX1_141/Y vdd INVX1
XINVX1_152 INVX1_152/A gnd NOR3X1_49/A vdd INVX1
XFILL_7_INVX1_138 gnd vdd FILL
XINVX1_163 NOR2X1_1/Y gnd INVX1_163/Y vdd INVX1
XFILL_7_INVX1_149 gnd vdd FILL
XINVX1_174 NAND2X1_6/B gnd INVX1_174/Y vdd INVX1
XINVX1_185 INVX1_185/A gnd NOR3X1_14/A vdd INVX1
XINVX1_196 INVX1_196/A gnd NOR3X1_41/A vdd INVX1
XFILL_22_NOR3X1_11 gnd vdd FILL
XFILL_15_MUX2X1_170 gnd vdd FILL
XFILL_22_NOR3X1_22 gnd vdd FILL
XFILL_22_NOR3X1_33 gnd vdd FILL
XFILL_15_MUX2X1_181 gnd vdd FILL
XFILL_72_DFFSR_200 gnd vdd FILL
XFILL_22_NOR3X1_44 gnd vdd FILL
XFILL_15_MUX2X1_192 gnd vdd FILL
XFILL_72_DFFSR_211 gnd vdd FILL
XFILL_72_DFFSR_222 gnd vdd FILL
XFILL_72_DFFSR_233 gnd vdd FILL
XFILL_72_DFFSR_244 gnd vdd FILL
XFILL_26_NOR3X1_10 gnd vdd FILL
XFILL_72_DFFSR_255 gnd vdd FILL
XFILL_72_DFFSR_266 gnd vdd FILL
XFILL_26_NOR3X1_21 gnd vdd FILL
XFILL_26_NOR3X1_32 gnd vdd FILL
XFILL_26_NOR3X1_43 gnd vdd FILL
XFILL_37_3_1 gnd vdd FILL
XFILL_76_DFFSR_210 gnd vdd FILL
XFILL_76_DFFSR_221 gnd vdd FILL
XFILL_76_DFFSR_232 gnd vdd FILL
XFILL_76_DFFSR_243 gnd vdd FILL
XFILL_1_NOR3X1_4 gnd vdd FILL
XFILL_76_DFFSR_254 gnd vdd FILL
XFILL_76_DFFSR_265 gnd vdd FILL
XFILL_31_CLKBUF1_6 gnd vdd FILL
XFILL_9_AOI21X1_17 gnd vdd FILL
XFILL_9_AOI21X1_28 gnd vdd FILL
XFILL_9_AOI21X1_39 gnd vdd FILL
XFILL_19_OAI22X1_19 gnd vdd FILL
XFILL_21_7_2 gnd vdd FILL
XFILL_35_CLKBUF1_5 gnd vdd FILL
XFILL_20_CLKBUF1_16 gnd vdd FILL
XFILL_20_2_1 gnd vdd FILL
XFILL_20_CLKBUF1_27 gnd vdd FILL
XFILL_20_CLKBUF1_38 gnd vdd FILL
XFILL_43_DFFSR_4 gnd vdd FILL
XFILL_6_BUFX2_9 gnd vdd FILL
XFILL_1_NOR2X1_105 gnd vdd FILL
XFILL_1_NOR2X1_116 gnd vdd FILL
XFILL_1_NOR2X1_127 gnd vdd FILL
XFILL_1_NOR2X1_138 gnd vdd FILL
XFILL_1_NOR2X1_149 gnd vdd FILL
XFILL_65_DFFSR_8 gnd vdd FILL
XFILL_8_BUFX4_17 gnd vdd FILL
XFILL_11_NAND2X1_20 gnd vdd FILL
XFILL_8_BUFX4_28 gnd vdd FILL
XFILL_11_NAND2X1_31 gnd vdd FILL
XFILL_11_NAND2X1_42 gnd vdd FILL
XFILL_11_NAND2X1_53 gnd vdd FILL
XFILL_1_OAI21X1_1 gnd vdd FILL
XFILL_8_BUFX4_39 gnd vdd FILL
XFILL_11_NAND2X1_64 gnd vdd FILL
XFILL_9_OAI22X1_14 gnd vdd FILL
XFILL_9_OAI22X1_25 gnd vdd FILL
XFILL_11_NAND2X1_75 gnd vdd FILL
XFILL_28_3_1 gnd vdd FILL
XFILL_3_3_1 gnd vdd FILL
XFILL_11_NAND2X1_86 gnd vdd FILL
XFILL_9_OAI22X1_36 gnd vdd FILL
XFILL_9_OAI22X1_47 gnd vdd FILL
XFILL_43_DFFSR_210 gnd vdd FILL
XFILL_43_DFFSR_221 gnd vdd FILL
XFILL_43_DFFSR_232 gnd vdd FILL
XFILL_43_DFFSR_243 gnd vdd FILL
XFILL_43_DFFSR_254 gnd vdd FILL
XFILL_43_DFFSR_265 gnd vdd FILL
XNAND3X1_105 DFFSR_79/Q BUFX4_58/Y AND2X2_5/Y gnd NAND3X1_106/C vdd NAND3X1
XFILL_2_NOR2X1_80 gnd vdd FILL
XNAND3X1_116 DFFSR_181/Q BUFX4_91/Y NOR2X1_30/Y gnd NAND3X1_118/A vdd NAND3X1
XFILL_2_NOR2X1_91 gnd vdd FILL
XNAND3X1_127 NAND2X1_72/Y NOR2X1_89/Y NOR3X1_32/Y gnd NOR2X1_91/B vdd NAND3X1
XFILL_8_NAND3X1_90 gnd vdd FILL
XFILL_5_BUFX4_3 gnd vdd FILL
XFILL_70_DFFSR_110 gnd vdd FILL
XFILL_6_NOR2X1_205 gnd vdd FILL
XFILL_47_DFFSR_220 gnd vdd FILL
XFILL_70_DFFSR_121 gnd vdd FILL
XFILL_70_DFFSR_132 gnd vdd FILL
XFILL_12_7_2 gnd vdd FILL
XFILL_47_DFFSR_231 gnd vdd FILL
XFILL_70_DFFSR_143 gnd vdd FILL
XFILL_70_DFFSR_154 gnd vdd FILL
XFILL_47_DFFSR_242 gnd vdd FILL
XFILL_47_DFFSR_253 gnd vdd FILL
XFILL_11_2_1 gnd vdd FILL
XFILL_15_AND2X2_5 gnd vdd FILL
XFILL_70_DFFSR_165 gnd vdd FILL
XFILL_47_DFFSR_264 gnd vdd FILL
XFILL_47_DFFSR_275 gnd vdd FILL
XFILL_70_DFFSR_176 gnd vdd FILL
XFILL_6_NOR2X1_90 gnd vdd FILL
XFILL_2_OAI21X1_16 gnd vdd FILL
XFILL_70_DFFSR_187 gnd vdd FILL
XFILL_2_OAI21X1_27 gnd vdd FILL
XFILL_70_DFFSR_198 gnd vdd FILL
XFILL_2_OAI21X1_38 gnd vdd FILL
XFILL_74_DFFSR_120 gnd vdd FILL
XFILL_2_OAI21X1_49 gnd vdd FILL
XFILL_74_DFFSR_131 gnd vdd FILL
XFILL_74_DFFSR_142 gnd vdd FILL
XFILL_74_DFFSR_153 gnd vdd FILL
XFILL_15_AOI21X1_20 gnd vdd FILL
XFILL_74_DFFSR_164 gnd vdd FILL
XFILL_15_AOI21X1_31 gnd vdd FILL
XFILL_15_AOI21X1_42 gnd vdd FILL
XFILL_74_DFFSR_175 gnd vdd FILL
XFILL_74_DFFSR_186 gnd vdd FILL
XFILL_15_AOI21X1_53 gnd vdd FILL
XFILL_74_DFFSR_197 gnd vdd FILL
XFILL_15_AOI21X1_64 gnd vdd FILL
XFILL_12_BUFX4_11 gnd vdd FILL
XFILL_12_BUFX4_22 gnd vdd FILL
XFILL_15_AOI21X1_75 gnd vdd FILL
XFILL_1_NAND2X1_70 gnd vdd FILL
XFILL_78_DFFSR_130 gnd vdd FILL
XFILL_1_NAND2X1_81 gnd vdd FILL
XFILL_4_INVX1_7 gnd vdd FILL
XFILL_12_BUFX4_33 gnd vdd FILL
XFILL_78_DFFSR_141 gnd vdd FILL
XFILL_78_DFFSR_152 gnd vdd FILL
XFILL_1_NAND2X1_92 gnd vdd FILL
XFILL_12_BUFX4_44 gnd vdd FILL
XFILL_78_DFFSR_163 gnd vdd FILL
XFILL_12_BUFX4_55 gnd vdd FILL
XFILL_78_DFFSR_174 gnd vdd FILL
XFILL_12_BUFX4_66 gnd vdd FILL
XFILL_12_BUFX4_77 gnd vdd FILL
XFILL_78_DFFSR_185 gnd vdd FILL
XFILL_12_BUFX4_88 gnd vdd FILL
XFILL_78_DFFSR_196 gnd vdd FILL
XFILL_12_BUFX4_99 gnd vdd FILL
XFILL_29_DFFSR_209 gnd vdd FILL
XFILL_56_DFFSR_109 gnd vdd FILL
XFILL_2_NAND2X1_2 gnd vdd FILL
XFILL_19_3_1 gnd vdd FILL
XFILL_62_6_2 gnd vdd FILL
XFILL_6_NAND2X1_1 gnd vdd FILL
XFILL_6_INVX1_12 gnd vdd FILL
XFILL_6_INVX1_23 gnd vdd FILL
XFILL_6_INVX1_34 gnd vdd FILL
XFILL_61_1_1 gnd vdd FILL
XFILL_18_MUX2X1_103 gnd vdd FILL
XFILL_8_INVX8_1 gnd vdd FILL
XFILL_10_DFFSR_210 gnd vdd FILL
XFILL_18_MUX2X1_114 gnd vdd FILL
XFILL_6_INVX1_45 gnd vdd FILL
XFILL_10_DFFSR_221 gnd vdd FILL
XFILL_7_AND2X2_4 gnd vdd FILL
XFILL_6_INVX1_56 gnd vdd FILL
XFILL_18_MUX2X1_125 gnd vdd FILL
XFILL_10_DFFSR_232 gnd vdd FILL
XFILL_20_5 gnd vdd FILL
XFILL_10_DFFSR_243 gnd vdd FILL
XFILL_6_INVX1_67 gnd vdd FILL
XFILL_18_MUX2X1_136 gnd vdd FILL
XFILL_10_DFFSR_254 gnd vdd FILL
XFILL_6_INVX1_78 gnd vdd FILL
XFILL_18_MUX2X1_147 gnd vdd FILL
XFILL_6_INVX1_89 gnd vdd FILL
XFILL_18_MUX2X1_158 gnd vdd FILL
XFILL_10_DFFSR_265 gnd vdd FILL
XFILL_5_AOI21X1_70 gnd vdd FILL
XFILL_18_MUX2X1_169 gnd vdd FILL
XFILL_5_AOI21X1_81 gnd vdd FILL
XFILL_13_4 gnd vdd FILL
XFILL_15_OAI22X1_50 gnd vdd FILL
XFILL_14_DFFSR_220 gnd vdd FILL
XFILL_14_DFFSR_231 gnd vdd FILL
XFILL_14_DFFSR_242 gnd vdd FILL
XDFFSR_103 DFFSR_103/Q DFFSR_73/CLK DFFSR_73/R vdd DFFSR_103/D gnd vdd DFFSR
XFILL_14_DFFSR_253 gnd vdd FILL
XFILL_25_DFFSR_1 gnd vdd FILL
XFILL_4_BUFX4_10 gnd vdd FILL
XDFFSR_114 INVX1_184/A DFFSR_64/CLK DFFSR_2/R vdd DFFSR_114/D gnd vdd DFFSR
XFILL_14_DFFSR_264 gnd vdd FILL
XFILL_14_DFFSR_275 gnd vdd FILL
XFILL_4_BUFX4_21 gnd vdd FILL
XFILL_82_DFFSR_2 gnd vdd FILL
XDFFSR_125 INVX1_178/A DFFSR_2/CLK BUFX4_50/Y vdd DFFSR_125/D gnd vdd DFFSR
XFILL_4_BUFX4_32 gnd vdd FILL
XDFFSR_136 INVX1_161/A CLKBUF1_1/Y DFFSR_58/R vdd DFFSR_136/D gnd vdd DFFSR
XFILL_4_BUFX4_43 gnd vdd FILL
XFILL_8_NOR2X1_180 gnd vdd FILL
XFILL_8_NOR2X1_191 gnd vdd FILL
XDFFSR_147 INVX1_158/A DFFSR_55/CLK DFFSR_91/R vdd DFFSR_147/D gnd vdd DFFSR
XDFFSR_158 NOR2X1_90/A CLKBUF1_1/Y DFFSR_89/R vdd DFFSR_158/D gnd vdd DFFSR
XFILL_41_DFFSR_120 gnd vdd FILL
XFILL_4_BUFX4_54 gnd vdd FILL
XFILL_41_DFFSR_131 gnd vdd FILL
XFILL_2_AOI21X1_7 gnd vdd FILL
XFILL_4_BUFX4_65 gnd vdd FILL
XDFFSR_169 INVX1_145/A DFFSR_56/CLK DFFSR_42/R vdd MUX2X1_68/Y gnd vdd DFFSR
XFILL_18_DFFSR_230 gnd vdd FILL
XFILL_41_DFFSR_142 gnd vdd FILL
XFILL_4_BUFX4_76 gnd vdd FILL
XFILL_41_DFFSR_153 gnd vdd FILL
XFILL_18_DFFSR_241 gnd vdd FILL
XFILL_4_BUFX4_87 gnd vdd FILL
XFILL_18_DFFSR_252 gnd vdd FILL
XFILL_4_BUFX4_98 gnd vdd FILL
XFILL_18_DFFSR_263 gnd vdd FILL
XFILL_41_DFFSR_164 gnd vdd FILL
XFILL_18_DFFSR_274 gnd vdd FILL
XFILL_41_DFFSR_175 gnd vdd FILL
XFILL_41_DFFSR_186 gnd vdd FILL
XFILL_41_DFFSR_197 gnd vdd FILL
XFILL_15_MUX2X1_19 gnd vdd FILL
XFILL_45_DFFSR_130 gnd vdd FILL
XFILL_6_AOI21X1_6 gnd vdd FILL
XFILL_45_DFFSR_141 gnd vdd FILL
XFILL_45_DFFSR_152 gnd vdd FILL
XFILL_45_DFFSR_163 gnd vdd FILL
XFILL_22_MUX2X1_8 gnd vdd FILL
XFILL_45_DFFSR_174 gnd vdd FILL
XFILL_19_MUX2X1_18 gnd vdd FILL
XFILL_45_DFFSR_185 gnd vdd FILL
XFILL_45_DFFSR_196 gnd vdd FILL
XFILL_8_MUX2X1_120 gnd vdd FILL
XFILL_19_MUX2X1_29 gnd vdd FILL
XFILL_8_MUX2X1_131 gnd vdd FILL
XFILL_47_DFFSR_5 gnd vdd FILL
XFILL_49_DFFSR_140 gnd vdd FILL
XFILL_8_MUX2X1_142 gnd vdd FILL
XFILL_8_MUX2X1_153 gnd vdd FILL
XNOR3X1_14 NOR3X1_14/A NOR3X1_49/B NOR3X1_6/B gnd NOR3X1_17/B vdd NOR3X1
XFILL_49_DFFSR_151 gnd vdd FILL
XFILL_11_AOI22X1_3 gnd vdd FILL
XFILL_49_DFFSR_162 gnd vdd FILL
XFILL_8_MUX2X1_164 gnd vdd FILL
XNOR3X1_25 NOR3X1_25/A NOR3X1_25/B NOR3X1_25/C gnd NOR3X1_25/Y vdd NOR3X1
XFILL_8_MUX2X1_175 gnd vdd FILL
XNOR3X1_36 INVX1_66/Y NOR3X1_39/C INVX2_2/Y gnd NOR3X1_38/B vdd NOR3X1
XFILL_49_DFFSR_173 gnd vdd FILL
XNOR3X1_47 NOR3X1_47/A NOR3X1_47/B NOR3X1_47/C gnd NOR3X1_47/Y vdd NOR3X1
XFILL_8_MUX2X1_186 gnd vdd FILL
XFILL_49_DFFSR_184 gnd vdd FILL
XFILL_49_DFFSR_195 gnd vdd FILL
XFILL_23_DFFSR_109 gnd vdd FILL
XFILL_53_6_2 gnd vdd FILL
XFILL_15_AOI22X1_2 gnd vdd FILL
XFILL_52_1_1 gnd vdd FILL
XFILL_5_MUX2X1_9 gnd vdd FILL
XFILL_27_DFFSR_108 gnd vdd FILL
XFILL_27_DFFSR_119 gnd vdd FILL
XFILL_10_NAND3X1_17 gnd vdd FILL
XFILL_19_AOI22X1_1 gnd vdd FILL
XFILL_10_NAND3X1_28 gnd vdd FILL
XFILL_10_NAND3X1_39 gnd vdd FILL
XFILL_69_DFFSR_9 gnd vdd FILL
XFILL_39_DFFSR_10 gnd vdd FILL
XFILL_39_DFFSR_21 gnd vdd FILL
XFILL_30_CLKBUF1_17 gnd vdd FILL
XFILL_30_CLKBUF1_28 gnd vdd FILL
XFILL_39_DFFSR_32 gnd vdd FILL
XFILL_39_DFFSR_43 gnd vdd FILL
XFILL_30_CLKBUF1_39 gnd vdd FILL
XFILL_39_DFFSR_54 gnd vdd FILL
XFILL_39_DFFSR_65 gnd vdd FILL
XFILL_39_DFFSR_76 gnd vdd FILL
XFILL_39_DFFSR_87 gnd vdd FILL
XFILL_39_DFFSR_98 gnd vdd FILL
XFILL_79_DFFSR_20 gnd vdd FILL
XFILL_79_DFFSR_31 gnd vdd FILL
XFILL_73_DFFSR_209 gnd vdd FILL
XFILL_79_DFFSR_42 gnd vdd FILL
XFILL_0_DFFSR_17 gnd vdd FILL
XFILL_79_DFFSR_53 gnd vdd FILL
XFILL_0_DFFSR_28 gnd vdd FILL
XFILL_10_NOR2X1_5 gnd vdd FILL
XFILL_79_DFFSR_64 gnd vdd FILL
XFILL_0_DFFSR_39 gnd vdd FILL
XFILL_79_DFFSR_75 gnd vdd FILL
XFILL_79_DFFSR_86 gnd vdd FILL
XFILL_27_NOR3X1_19 gnd vdd FILL
XFILL_79_DFFSR_97 gnd vdd FILL
XFILL_9_BUFX4_4 gnd vdd FILL
XFILL_77_DFFSR_208 gnd vdd FILL
XFILL_2_INVX1_60 gnd vdd FILL
XFILL_12_DFFSR_130 gnd vdd FILL
XFILL_77_DFFSR_219 gnd vdd FILL
XFILL_2_INVX1_71 gnd vdd FILL
XFILL_12_DFFSR_141 gnd vdd FILL
XFILL_12_DFFSR_152 gnd vdd FILL
XFILL_2_INVX1_82 gnd vdd FILL
XFILL_2_INVX1_93 gnd vdd FILL
XFILL_48_DFFSR_30 gnd vdd FILL
XFILL_12_DFFSR_163 gnd vdd FILL
XFILL_48_DFFSR_41 gnd vdd FILL
XFILL_19_NOR3X1_5 gnd vdd FILL
XFILL_12_DFFSR_174 gnd vdd FILL
XFILL_1_CLKBUF1_6 gnd vdd FILL
XFILL_48_DFFSR_52 gnd vdd FILL
XFILL_12_DFFSR_185 gnd vdd FILL
XFILL_48_DFFSR_63 gnd vdd FILL
XFILL_12_DFFSR_196 gnd vdd FILL
XFILL_48_DFFSR_74 gnd vdd FILL
XFILL_0_NAND3X1_12 gnd vdd FILL
XFILL_48_DFFSR_85 gnd vdd FILL
XFILL_0_NAND3X1_23 gnd vdd FILL
XFILL_48_DFFSR_96 gnd vdd FILL
XFILL_16_DFFSR_140 gnd vdd FILL
XFILL_0_NAND3X1_34 gnd vdd FILL
XFILL_16_DFFSR_151 gnd vdd FILL
XFILL_0_NAND3X1_45 gnd vdd FILL
XFILL_16_DFFSR_162 gnd vdd FILL
XFILL_0_NAND3X1_56 gnd vdd FILL
XFILL_4_NAND2X1_14 gnd vdd FILL
XFILL_16_DFFSR_173 gnd vdd FILL
XFILL_0_NAND3X1_67 gnd vdd FILL
XFILL_4_NAND2X1_25 gnd vdd FILL
XFILL_5_CLKBUF1_5 gnd vdd FILL
XFILL_16_DFFSR_184 gnd vdd FILL
XFILL_0_NAND3X1_78 gnd vdd FILL
XFILL_4_NAND2X1_36 gnd vdd FILL
XFILL_44_6_2 gnd vdd FILL
XFILL_0_NAND3X1_89 gnd vdd FILL
XFILL_16_DFFSR_195 gnd vdd FILL
XFILL_4_NAND2X1_47 gnd vdd FILL
XFILL_17_DFFSR_40 gnd vdd FILL
XFILL_4_NAND2X1_58 gnd vdd FILL
XFILL_0_BUFX4_80 gnd vdd FILL
XFILL_17_DFFSR_51 gnd vdd FILL
XFILL_43_1_1 gnd vdd FILL
XFILL_4_NAND2X1_69 gnd vdd FILL
XFILL_0_BUFX4_91 gnd vdd FILL
XFILL_17_DFFSR_62 gnd vdd FILL
XFILL_1_BUFX4_100 gnd vdd FILL
XFILL_17_DFFSR_73 gnd vdd FILL
XFILL_17_DFFSR_84 gnd vdd FILL
XFILL_17_DFFSR_95 gnd vdd FILL
XFILL_9_CLKBUF1_4 gnd vdd FILL
XFILL_12_NOR3X1_30 gnd vdd FILL
XFILL_12_NOR3X1_41 gnd vdd FILL
XFILL_28_NOR3X1_3 gnd vdd FILL
XFILL_12_NOR3X1_52 gnd vdd FILL
XFILL_57_DFFSR_50 gnd vdd FILL
XFILL_57_DFFSR_61 gnd vdd FILL
XFILL_62_DFFSR_230 gnd vdd FILL
XFILL_57_DFFSR_72 gnd vdd FILL
XFILL_57_DFFSR_83 gnd vdd FILL
XFILL_62_DFFSR_241 gnd vdd FILL
XFILL_57_DFFSR_94 gnd vdd FILL
XFILL_62_DFFSR_252 gnd vdd FILL
XFILL_62_DFFSR_263 gnd vdd FILL
XFILL_62_DFFSR_274 gnd vdd FILL
XFILL_16_NOR3X1_40 gnd vdd FILL
XFILL_16_NOR3X1_51 gnd vdd FILL
XFILL_2_NOR2X1_4 gnd vdd FILL
XFILL_10_NOR2X1_107 gnd vdd FILL
XFILL_10_NOR2X1_118 gnd vdd FILL
XFILL_66_DFFSR_240 gnd vdd FILL
XFILL_10_NOR2X1_129 gnd vdd FILL
XFILL_66_DFFSR_251 gnd vdd FILL
XFILL_66_DFFSR_262 gnd vdd FILL
XFILL_26_DFFSR_60 gnd vdd FILL
XFILL_21_CLKBUF1_3 gnd vdd FILL
XFILL_66_DFFSR_273 gnd vdd FILL
XFILL_26_DFFSR_71 gnd vdd FILL
XFILL_26_DFFSR_82 gnd vdd FILL
XFILL_26_DFFSR_93 gnd vdd FILL
XFILL_40_DFFSR_209 gnd vdd FILL
XFILL_8_AOI21X1_14 gnd vdd FILL
XFILL_8_AOI21X1_25 gnd vdd FILL
XFILL_8_AOI21X1_36 gnd vdd FILL
XFILL_1_MUX2X1_2 gnd vdd FILL
XFILL_8_AOI21X1_47 gnd vdd FILL
XFILL_18_OAI22X1_16 gnd vdd FILL
XFILL_8_AOI21X1_58 gnd vdd FILL
XFILL_8_AOI21X1_69 gnd vdd FILL
XFILL_66_DFFSR_70 gnd vdd FILL
XFILL_25_CLKBUF1_2 gnd vdd FILL
XFILL_18_OAI22X1_27 gnd vdd FILL
XFILL_66_DFFSR_81 gnd vdd FILL
XFILL_18_OAI22X1_38 gnd vdd FILL
XFILL_3_NOR2X1_12 gnd vdd FILL
XFILL_66_DFFSR_92 gnd vdd FILL
XFILL_44_DFFSR_208 gnd vdd FILL
XFILL_3_NOR2X1_23 gnd vdd FILL
XFILL_18_OAI22X1_49 gnd vdd FILL
XFILL_44_DFFSR_219 gnd vdd FILL
XFILL_6_OAI21X1_9 gnd vdd FILL
XFILL_3_NOR2X1_34 gnd vdd FILL
XFILL_3_NOR2X1_45 gnd vdd FILL
XFILL_3_NOR2X1_56 gnd vdd FILL
XFILL_29_DFFSR_2 gnd vdd FILL
XFILL_3_NOR2X1_67 gnd vdd FILL
XFILL_86_DFFSR_3 gnd vdd FILL
XFILL_29_CLKBUF1_1 gnd vdd FILL
XNAND3X1_80 DFFSR_16/Q NAND3X1_7/B NOR2X1_36/Y gnd NAND3X1_82/B vdd NAND3X1
XFILL_2_CLKBUF1_17 gnd vdd FILL
XFILL_2_CLKBUF1_28 gnd vdd FILL
XNAND3X1_91 INVX1_161/A BUFX4_90/Y NOR3X1_51/Y gnd OAI21X1_11/C vdd NAND3X1
XFILL_3_NOR2X1_78 gnd vdd FILL
XFILL_9_DFFSR_50 gnd vdd FILL
XFILL_3_NOR2X1_89 gnd vdd FILL
XFILL_9_DFFSR_61 gnd vdd FILL
XFILL_2_CLKBUF1_39 gnd vdd FILL
XFILL_71_DFFSR_108 gnd vdd FILL
XFILL_7_NOR2X1_11 gnd vdd FILL
XFILL_9_DFFSR_72 gnd vdd FILL
XFILL_48_DFFSR_207 gnd vdd FILL
XFILL_7_NOR2X1_22 gnd vdd FILL
XFILL_9_DFFSR_83 gnd vdd FILL
XFILL_71_DFFSR_119 gnd vdd FILL
XFILL_48_DFFSR_218 gnd vdd FILL
XFILL_9_DFFSR_94 gnd vdd FILL
XFILL_7_NOR2X1_33 gnd vdd FILL
XFILL_48_DFFSR_229 gnd vdd FILL
XFILL_35_DFFSR_80 gnd vdd FILL
XFILL_35_6_2 gnd vdd FILL
XFILL_7_NOR2X1_44 gnd vdd FILL
XFILL_7_NOR2X1_55 gnd vdd FILL
XFILL_11_OAI22X1_6 gnd vdd FILL
XFILL_35_DFFSR_91 gnd vdd FILL
XNOR2X1_80 INVX1_38/Y NOR2X1_80/B gnd NOR3X1_30/B vdd NOR2X1
XFILL_7_NOR2X1_66 gnd vdd FILL
XFILL_7_NOR2X1_77 gnd vdd FILL
XFILL_34_1_1 gnd vdd FILL
XNOR2X1_91 NOR2X1_91/A NOR2X1_91/B gnd NOR2X1_91/Y vdd NOR2X1
XFILL_7_NOR2X1_88 gnd vdd FILL
XFILL_75_DFFSR_107 gnd vdd FILL
XFILL_0_NOR2X1_102 gnd vdd FILL
XFILL_7_NOR2X1_99 gnd vdd FILL
XFILL_0_NOR2X1_113 gnd vdd FILL
XFILL_75_DFFSR_118 gnd vdd FILL
XFILL_11_OAI21X1_18 gnd vdd FILL
XFILL_0_NOR2X1_124 gnd vdd FILL
XFILL_11_OAI21X1_29 gnd vdd FILL
XFILL_75_DFFSR_129 gnd vdd FILL
XFILL_0_NOR2X1_135 gnd vdd FILL
XFILL_75_DFFSR_90 gnd vdd FILL
XFILL_0_NOR2X1_146 gnd vdd FILL
XFILL_15_OAI22X1_5 gnd vdd FILL
XFILL_0_NOR2X1_157 gnd vdd FILL
XFILL_13_DFFSR_8 gnd vdd FILL
XFILL_11_1 gnd vdd FILL
XFILL_0_NOR2X1_168 gnd vdd FILL
XFILL_70_DFFSR_9 gnd vdd FILL
XFILL_0_NOR2X1_179 gnd vdd FILL
XFILL_79_DFFSR_106 gnd vdd FILL
XFILL_79_DFFSR_117 gnd vdd FILL
XFILL_10_NAND2X1_50 gnd vdd FILL
XFILL_79_DFFSR_128 gnd vdd FILL
XFILL_10_NAND2X1_61 gnd vdd FILL
XFILL_79_DFFSR_139 gnd vdd FILL
XFILL_19_OAI22X1_4 gnd vdd FILL
XFILL_10_NAND2X1_72 gnd vdd FILL
XFILL_8_OAI22X1_11 gnd vdd FILL
XFILL_8_OAI22X1_22 gnd vdd FILL
XFILL_10_NAND2X1_83 gnd vdd FILL
XFILL_8_OAI22X1_33 gnd vdd FILL
XFILL_10_NAND2X1_94 gnd vdd FILL
XFILL_8_OAI22X1_44 gnd vdd FILL
XBUFX2_7 BUFX2_7/A gnd addr[3] vdd BUFX2
XFILL_24_10 gnd vdd FILL
XFILL_33_DFFSR_240 gnd vdd FILL
XFILL_33_DFFSR_251 gnd vdd FILL
XFILL_33_DFFSR_262 gnd vdd FILL
XFILL_33_DFFSR_273 gnd vdd FILL
XFILL_0_MUX2X1_108 gnd vdd FILL
XFILL_0_MUX2X1_119 gnd vdd FILL
XFILL_5_NOR2X1_202 gnd vdd FILL
XFILL_60_DFFSR_140 gnd vdd FILL
XFILL_60_DFFSR_151 gnd vdd FILL
XFILL_60_DFFSR_162 gnd vdd FILL
XFILL_37_DFFSR_250 gnd vdd FILL
XNAND2X1_2 INVX4_1/A INVX1_8/A gnd NAND2X1_2/Y vdd NAND2X1
XFILL_37_DFFSR_261 gnd vdd FILL
XFILL_1_OAI21X1_13 gnd vdd FILL
XFILL_37_DFFSR_272 gnd vdd FILL
XFILL_60_DFFSR_173 gnd vdd FILL
XFILL_60_DFFSR_184 gnd vdd FILL
XFILL_1_OAI21X1_24 gnd vdd FILL
XFILL_3_MUX2X1_30 gnd vdd FILL
XFILL_60_DFFSR_195 gnd vdd FILL
XFILL_19_CLKBUF1_20 gnd vdd FILL
XFILL_11_DFFSR_208 gnd vdd FILL
XFILL_1_OAI21X1_35 gnd vdd FILL
XFILL_3_MUX2X1_41 gnd vdd FILL
XFILL_11_DFFSR_219 gnd vdd FILL
XFILL_3_MUX2X1_52 gnd vdd FILL
XFILL_1_OAI21X1_46 gnd vdd FILL
XFILL_19_CLKBUF1_31 gnd vdd FILL
XFILL_3_MUX2X1_63 gnd vdd FILL
XFILL_19_CLKBUF1_42 gnd vdd FILL
XFILL_3_MUX2X1_74 gnd vdd FILL
XFILL_64_DFFSR_150 gnd vdd FILL
XFILL_64_DFFSR_161 gnd vdd FILL
XFILL_3_MUX2X1_85 gnd vdd FILL
XFILL_3_MUX2X1_96 gnd vdd FILL
XFILL_64_DFFSR_172 gnd vdd FILL
XFILL_14_AOI21X1_50 gnd vdd FILL
XFILL_64_DFFSR_183 gnd vdd FILL
XFILL_26_6_2 gnd vdd FILL
XFILL_1_6_2 gnd vdd FILL
XFILL_64_DFFSR_194 gnd vdd FILL
XFILL_14_AOI21X1_61 gnd vdd FILL
XFILL_15_DFFSR_207 gnd vdd FILL
XFILL_14_AOI21X1_72 gnd vdd FILL
XFILL_7_MUX2X1_40 gnd vdd FILL
XFILL_7_MUX2X1_51 gnd vdd FILL
XFILL_12_NAND3X1_7 gnd vdd FILL
XFILL_15_DFFSR_218 gnd vdd FILL
XFILL_25_1_1 gnd vdd FILL
XFILL_7_MUX2X1_62 gnd vdd FILL
XFILL_0_1_1 gnd vdd FILL
XFILL_15_DFFSR_229 gnd vdd FILL
XFILL_7_MUX2X1_73 gnd vdd FILL
XFILL_68_DFFSR_160 gnd vdd FILL
XFILL_7_MUX2X1_84 gnd vdd FILL
XNOR2X1_170 NOR2X1_20/A NAND2X1_3/Y gnd MUX2X1_3/S vdd NOR2X1
XFILL_7_MUX2X1_95 gnd vdd FILL
XFILL_68_DFFSR_171 gnd vdd FILL
XNOR2X1_181 DFFSR_31/Q NOR2X1_181/B gnd NOR2X1_181/Y vdd NOR2X1
XFILL_68_DFFSR_182 gnd vdd FILL
XNOR2X1_192 DFFSR_15/Q NOR2X1_195/B gnd NOR2X1_192/Y vdd NOR2X1
XFILL_42_DFFSR_107 gnd vdd FILL
XFILL_68_DFFSR_193 gnd vdd FILL
XFILL_19_DFFSR_206 gnd vdd FILL
XFILL_19_DFFSR_217 gnd vdd FILL
XFILL_42_DFFSR_118 gnd vdd FILL
XFILL_19_DFFSR_228 gnd vdd FILL
XFILL_42_DFFSR_129 gnd vdd FILL
XFILL_19_DFFSR_239 gnd vdd FILL
XFILL_46_DFFSR_106 gnd vdd FILL
XFILL_46_DFFSR_117 gnd vdd FILL
XAOI21X1_7 BUFX4_99/Y AOI21X1_7/B AOI21X1_7/C gnd DFFSR_142/D vdd AOI21X1
XFILL_46_DFFSR_128 gnd vdd FILL
XFILL_46_DFFSR_139 gnd vdd FILL
XMUX2X1_110 NOR2X1_62/A BUFX4_67/Y NAND2X1_23/Y gnd DFFSR_153/D vdd MUX2X1
XMUX2X1_121 INVX1_164/Y MUX2X1_2/A NAND2X1_78/Y gnd DFFSR_138/D vdd MUX2X1
XMUX2X1_132 INVX1_176/Y BUFX4_66/Y NAND2X1_2/Y gnd DFFSR_122/D vdd MUX2X1
XFILL_17_MUX2X1_100 gnd vdd FILL
XMUX2X1_143 INVX1_187/Y BUFX4_93/Y NAND3X1_1/Y gnd DFFSR_116/D vdd MUX2X1
XFILL_17_MUX2X1_111 gnd vdd FILL
XMUX2X1_154 MUX2X1_1/A INVX1_198/Y NOR2X1_155/Y gnd DFFSR_91/D vdd MUX2X1
XMUX2X1_165 BUFX4_98/Y INVX1_210/Y NOR2X1_162/Y gnd DFFSR_80/D vdd MUX2X1
XFILL_17_MUX2X1_122 gnd vdd FILL
XFILL_23_MUX2X1_60 gnd vdd FILL
XMUX2X1_176 BUFX4_67/Y OAI22X1_9/A NOR2X1_166/Y gnd DFFSR_64/D vdd MUX2X1
XFILL_23_MUX2X1_71 gnd vdd FILL
XFILL_9_7_2 gnd vdd FILL
XFILL_17_MUX2X1_133 gnd vdd FILL
XFILL_17_MUX2X1_144 gnd vdd FILL
XMUX2X1_187 BUFX4_99/Y INVX1_6/Y NOR2X1_168/Y gnd DFFSR_58/D vdd MUX2X1
XFILL_17_MUX2X1_155 gnd vdd FILL
XFILL_23_MUX2X1_82 gnd vdd FILL
XFILL_9_BUFX2_1 gnd vdd FILL
XFILL_23_MUX2X1_93 gnd vdd FILL
XFILL_8_2_1 gnd vdd FILL
XFILL_17_MUX2X1_166 gnd vdd FILL
XFILL_17_MUX2X1_177 gnd vdd FILL
XFILL_17_MUX2X1_188 gnd vdd FILL
XINVX1_50 INVX1_50/A gnd INVX1_50/Y vdd INVX1
XFILL_30_DFFSR_2 gnd vdd FILL
XINVX1_61 INVX1_61/A gnd INVX1_61/Y vdd INVX1
XINVX1_72 INVX1_72/A gnd INVX1_72/Y vdd INVX1
XINVX1_83 INVX1_83/A gnd INVX1_83/Y vdd INVX1
XINVX1_94 INVX1_94/A gnd INVX1_94/Y vdd INVX1
XFILL_3_INVX1_16 gnd vdd FILL
XFILL_3_INVX1_27 gnd vdd FILL
XFILL_3_INVX1_38 gnd vdd FILL
XFILL_31_DFFSR_150 gnd vdd FILL
XFILL_17_6_2 gnd vdd FILL
XFILL_31_DFFSR_161 gnd vdd FILL
XFILL_3_INVX1_49 gnd vdd FILL
XFILL_4_AND2X2_8 gnd vdd FILL
XFILL_31_DFFSR_172 gnd vdd FILL
XFILL_16_1_1 gnd vdd FILL
XFILL_31_DFFSR_183 gnd vdd FILL
XFILL_49_DFFSR_19 gnd vdd FILL
XFILL_31_DFFSR_194 gnd vdd FILL
XFILL_35_DFFSR_160 gnd vdd FILL
XFILL_35_DFFSR_171 gnd vdd FILL
XFILL_35_DFFSR_182 gnd vdd FILL
XFILL_35_DFFSR_193 gnd vdd FILL
XFILL_1_BUFX4_14 gnd vdd FILL
XFILL_52_DFFSR_6 gnd vdd FILL
XFILL_1_BUFX4_25 gnd vdd FILL
XFILL_1_BUFX4_36 gnd vdd FILL
XFILL_1_BUFX4_47 gnd vdd FILL
XFILL_7_MUX2X1_150 gnd vdd FILL
XFILL_18_DFFSR_18 gnd vdd FILL
XFILL_7_MUX2X1_161 gnd vdd FILL
XFILL_18_DFFSR_29 gnd vdd FILL
XFILL_1_BUFX4_58 gnd vdd FILL
XFILL_39_DFFSR_170 gnd vdd FILL
XFILL_1_BUFX4_69 gnd vdd FILL
XFILL_7_MUX2X1_172 gnd vdd FILL
XFILL_7_MUX2X1_183 gnd vdd FILL
XFILL_39_DFFSR_181 gnd vdd FILL
XFILL_7_MUX2X1_194 gnd vdd FILL
XFILL_13_DFFSR_106 gnd vdd FILL
XFILL_39_DFFSR_192 gnd vdd FILL
XFILL_13_DFFSR_117 gnd vdd FILL
XFILL_31_NOR3X1_50 gnd vdd FILL
XFILL_13_DFFSR_128 gnd vdd FILL
XFILL_13_DFFSR_139 gnd vdd FILL
XFILL_58_DFFSR_17 gnd vdd FILL
XNOR2X1_5 NOR2X1_5/A NOR2X1_6/B gnd NOR2X1_5/Y vdd NOR2X1
XFILL_58_DFFSR_28 gnd vdd FILL
XFILL_58_DFFSR_39 gnd vdd FILL
XFILL_81_DFFSR_250 gnd vdd FILL
XFILL_81_DFFSR_261 gnd vdd FILL
XFILL_17_DFFSR_105 gnd vdd FILL
XFILL_81_DFFSR_272 gnd vdd FILL
XFILL_17_DFFSR_116 gnd vdd FILL
XFILL_17_DFFSR_127 gnd vdd FILL
XFILL_17_DFFSR_138 gnd vdd FILL
XFILL_17_DFFSR_149 gnd vdd FILL
XFILL_12_AOI21X1_1 gnd vdd FILL
XFILL_17_DFFSR_9 gnd vdd FILL
XFILL_85_DFFSR_260 gnd vdd FILL
XFILL_85_DFFSR_271 gnd vdd FILL
XFILL_27_DFFSR_16 gnd vdd FILL
XFILL_66_2 gnd vdd FILL
XFILL_27_DFFSR_27 gnd vdd FILL
XFILL_27_DFFSR_38 gnd vdd FILL
XFILL_27_DFFSR_49 gnd vdd FILL
XFILL_66_0_1 gnd vdd FILL
XFILL_59_1 gnd vdd FILL
XFILL_13_NOR3X1_17 gnd vdd FILL
XFILL_67_DFFSR_15 gnd vdd FILL
XFILL_13_NOR3X1_28 gnd vdd FILL
XFILL_67_DFFSR_26 gnd vdd FILL
XFILL_13_NOR3X1_39 gnd vdd FILL
XFILL_67_DFFSR_37 gnd vdd FILL
XFILL_63_DFFSR_206 gnd vdd FILL
XFILL_67_DFFSR_48 gnd vdd FILL
XFILL_63_DFFSR_217 gnd vdd FILL
XFILL_67_DFFSR_59 gnd vdd FILL
XFILL_63_DFFSR_228 gnd vdd FILL
XFILL_63_DFFSR_239 gnd vdd FILL
XFILL_17_NOR3X1_16 gnd vdd FILL
XFILL_17_NOR3X1_27 gnd vdd FILL
XFILL_50_4_2 gnd vdd FILL
XFILL_17_NOR3X1_38 gnd vdd FILL
XFILL_17_NOR3X1_49 gnd vdd FILL
XFILL_67_DFFSR_205 gnd vdd FILL
XFILL_67_DFFSR_216 gnd vdd FILL
XFILL_36_DFFSR_14 gnd vdd FILL
XFILL_67_DFFSR_227 gnd vdd FILL
XFILL_36_DFFSR_25 gnd vdd FILL
XFILL_67_DFFSR_238 gnd vdd FILL
XFILL_36_DFFSR_36 gnd vdd FILL
XFILL_67_DFFSR_249 gnd vdd FILL
XFILL_36_DFFSR_47 gnd vdd FILL
XFILL_36_DFFSR_58 gnd vdd FILL
XFILL_36_DFFSR_69 gnd vdd FILL
XAOI21X1_15 BUFX4_78/Y NOR2X1_153/B NOR2X1_151/Y gnd DFFSR_100/D vdd AOI21X1
XAOI21X1_26 MUX2X1_6/B NOR2X1_181/B NOR2X1_180/Y gnd DFFSR_30/D vdd AOI21X1
XFILL_76_DFFSR_13 gnd vdd FILL
XFILL_76_DFFSR_24 gnd vdd FILL
XAOI21X1_37 BUFX4_78/Y NOR2X1_195/B NOR2X1_194/Y gnd DFFSR_17/D vdd AOI21X1
XFILL_76_DFFSR_35 gnd vdd FILL
XAOI21X1_48 BUFX4_71/Y NOR2X1_6/B NOR2X1_5/Y gnd DFFSR_273/D vdd AOI21X1
XAOI21X1_59 BUFX4_75/Y NOR2X1_26/B NOR2X1_26/Y gnd DFFSR_207/D vdd AOI21X1
XFILL_3_NAND2X1_11 gnd vdd FILL
XFILL_76_DFFSR_46 gnd vdd FILL
XFILL_19_MUX2X1_3 gnd vdd FILL
XFILL_76_DFFSR_57 gnd vdd FILL
XFILL_3_NAND2X1_22 gnd vdd FILL
XFILL_76_DFFSR_68 gnd vdd FILL
XFILL_3_NAND2X1_33 gnd vdd FILL
XFILL_76_DFFSR_79 gnd vdd FILL
XFILL_3_NAND2X1_44 gnd vdd FILL
XFILL_3_NAND2X1_55 gnd vdd FILL
XFILL_3_NAND2X1_66 gnd vdd FILL
XFILL_11_BUFX4_9 gnd vdd FILL
XFILL_3_NAND2X1_77 gnd vdd FILL
XFILL_0_AND2X2_1 gnd vdd FILL
XFILL_3_NAND2X1_88 gnd vdd FILL
XFILL_45_DFFSR_12 gnd vdd FILL
XFILL_45_DFFSR_23 gnd vdd FILL
XFILL_45_DFFSR_34 gnd vdd FILL
XFILL_11_CLKBUF1_19 gnd vdd FILL
XFILL_16_NOR3X1_9 gnd vdd FILL
XFILL_45_DFFSR_45 gnd vdd FILL
XFILL_45_DFFSR_56 gnd vdd FILL
XFILL_45_DFFSR_67 gnd vdd FILL
XFILL_45_DFFSR_78 gnd vdd FILL
XFILL_45_DFFSR_89 gnd vdd FILL
XFILL_58_5_2 gnd vdd FILL
XFILL_85_DFFSR_11 gnd vdd FILL
XFILL_57_0_1 gnd vdd FILL
XFILL_85_DFFSR_22 gnd vdd FILL
XFILL_52_DFFSR_260 gnd vdd FILL
XFILL_52_DFFSR_271 gnd vdd FILL
XFILL_85_DFFSR_33 gnd vdd FILL
XFILL_85_DFFSR_44 gnd vdd FILL
XFILL_85_DFFSR_55 gnd vdd FILL
XFILL_29_CLKBUF1_10 gnd vdd FILL
XFILL_29_CLKBUF1_21 gnd vdd FILL
XFILL_14_DFFSR_11 gnd vdd FILL
XFILL_29_CLKBUF1_32 gnd vdd FILL
XFILL_14_DFFSR_22 gnd vdd FILL
XFILL_85_DFFSR_66 gnd vdd FILL
XFILL_85_DFFSR_77 gnd vdd FILL
XFILL_14_DFFSR_33 gnd vdd FILL
XFILL_85_DFFSR_88 gnd vdd FILL
XFILL_14_DFFSR_44 gnd vdd FILL
XFILL_14_DFFSR_55 gnd vdd FILL
XFILL_85_DFFSR_99 gnd vdd FILL
XFILL_14_DFFSR_66 gnd vdd FILL
XFILL_14_DFFSR_77 gnd vdd FILL
XFILL_56_DFFSR_270 gnd vdd FILL
XFILL_14_DFFSR_88 gnd vdd FILL
XFILL_14_DFFSR_99 gnd vdd FILL
XFILL_54_DFFSR_10 gnd vdd FILL
XFILL_30_DFFSR_206 gnd vdd FILL
XFILL_7_AOI21X1_11 gnd vdd FILL
XFILL_54_DFFSR_21 gnd vdd FILL
XFILL_30_DFFSR_217 gnd vdd FILL
XOAI22X1_12 INVX1_54/Y OAI22X1_33/B INVX1_59/Y OAI22X1_33/D gnd NOR2X1_33/B vdd OAI22X1
XFILL_7_AOI21X1_22 gnd vdd FILL
XOAI22X1_23 INVX1_45/Y OAI22X1_32/B INVX1_50/Y OAI22X1_32/D gnd NOR2X1_33/A vdd OAI22X1
XFILL_30_DFFSR_228 gnd vdd FILL
XFILL_54_DFFSR_32 gnd vdd FILL
XFILL_54_DFFSR_43 gnd vdd FILL
XFILL_7_AOI21X1_33 gnd vdd FILL
XOAI22X1_34 MUX2X1_4/A OAI21X1_8/B INVX1_28/Y OAI22X1_36/B gnd NOR2X1_39/A vdd OAI22X1
XFILL_25_NOR3X1_7 gnd vdd FILL
XFILL_7_AOI21X1_44 gnd vdd FILL
XFILL_41_4_2 gnd vdd FILL
XFILL_30_DFFSR_239 gnd vdd FILL
XFILL_54_DFFSR_54 gnd vdd FILL
XFILL_54_DFFSR_65 gnd vdd FILL
XOAI22X1_45 INVX1_220/Y OAI22X1_9/B INVX1_224/Y OAI22X1_9/D gnd NOR2X1_48/B vdd OAI22X1
XFILL_83_DFFSR_170 gnd vdd FILL
XFILL_7_AOI21X1_55 gnd vdd FILL
XFILL_17_OAI22X1_13 gnd vdd FILL
XFILL_54_DFFSR_76 gnd vdd FILL
XFILL_7_AOI21X1_66 gnd vdd FILL
XFILL_17_OAI22X1_24 gnd vdd FILL
XFILL_54_DFFSR_87 gnd vdd FILL
XFILL_7_AOI21X1_77 gnd vdd FILL
XFILL_83_DFFSR_181 gnd vdd FILL
XFILL_54_DFFSR_98 gnd vdd FILL
XFILL_17_OAI22X1_35 gnd vdd FILL
XFILL_83_DFFSR_192 gnd vdd FILL
XFILL_34_DFFSR_205 gnd vdd FILL
XFILL_17_OAI22X1_46 gnd vdd FILL
XFILL_34_DFFSR_216 gnd vdd FILL
XFILL_34_DFFSR_227 gnd vdd FILL
XFILL_3_DFFSR_240 gnd vdd FILL
XFILL_34_DFFSR_3 gnd vdd FILL
XFILL_34_DFFSR_238 gnd vdd FILL
XFILL_3_DFFSR_251 gnd vdd FILL
XFILL_34_DFFSR_249 gnd vdd FILL
XFILL_3_DFFSR_262 gnd vdd FILL
XFILL_23_DFFSR_20 gnd vdd FILL
XFILL_3_DFFSR_273 gnd vdd FILL
XFILL_1_CLKBUF1_14 gnd vdd FILL
XFILL_1_CLKBUF1_25 gnd vdd FILL
XFILL_87_DFFSR_180 gnd vdd FILL
XFILL_0_MUX2X1_18 gnd vdd FILL
XFILL_23_DFFSR_31 gnd vdd FILL
XFILL_1_CLKBUF1_36 gnd vdd FILL
XFILL_23_DFFSR_42 gnd vdd FILL
XFILL_61_DFFSR_105 gnd vdd FILL
XFILL_0_MUX2X1_29 gnd vdd FILL
XFILL_23_DFFSR_53 gnd vdd FILL
XFILL_87_DFFSR_191 gnd vdd FILL
XFILL_61_DFFSR_116 gnd vdd FILL
XFILL_23_DFFSR_64 gnd vdd FILL
XFILL_38_DFFSR_204 gnd vdd FILL
XFILL_38_DFFSR_215 gnd vdd FILL
XFILL_23_DFFSR_75 gnd vdd FILL
XFILL_61_DFFSR_127 gnd vdd FILL
XFILL_38_DFFSR_226 gnd vdd FILL
XFILL_61_DFFSR_138 gnd vdd FILL
XFILL_23_DFFSR_86 gnd vdd FILL
XFILL_38_DFFSR_237 gnd vdd FILL
XFILL_7_DFFSR_250 gnd vdd FILL
XFILL_61_DFFSR_149 gnd vdd FILL
XFILL_23_DFFSR_97 gnd vdd FILL
XFILL_8_NOR3X1_8 gnd vdd FILL
XFILL_38_DFFSR_248 gnd vdd FILL
XFILL_7_DFFSR_261 gnd vdd FILL
XFILL_7_DFFSR_272 gnd vdd FILL
XFILL_63_DFFSR_30 gnd vdd FILL
XFILL_38_DFFSR_259 gnd vdd FILL
XFILL_4_MUX2X1_17 gnd vdd FILL
XFILL_63_DFFSR_41 gnd vdd FILL
XFILL_65_DFFSR_104 gnd vdd FILL
XFILL_63_DFFSR_52 gnd vdd FILL
XFILL_4_MUX2X1_28 gnd vdd FILL
XFILL_63_DFFSR_63 gnd vdd FILL
XFILL_4_MUX2X1_39 gnd vdd FILL
XFILL_65_DFFSR_115 gnd vdd FILL
XFILL_10_OAI21X1_15 gnd vdd FILL
XFILL_63_DFFSR_74 gnd vdd FILL
XFILL_10_OAI21X1_26 gnd vdd FILL
XFILL_63_DFFSR_85 gnd vdd FILL
XFILL_65_DFFSR_126 gnd vdd FILL
XFILL_65_DFFSR_137 gnd vdd FILL
XFILL_10_OAI21X1_37 gnd vdd FILL
XFILL_65_DFFSR_148 gnd vdd FILL
XFILL_63_DFFSR_96 gnd vdd FILL
XFILL_10_OAI21X1_48 gnd vdd FILL
XFILL_65_DFFSR_159 gnd vdd FILL
XFILL_6_DFFSR_10 gnd vdd FILL
XFILL_6_DFFSR_21 gnd vdd FILL
XFILL_8_MUX2X1_16 gnd vdd FILL
XFILL_8_MUX2X1_27 gnd vdd FILL
XFILL_69_DFFSR_103 gnd vdd FILL
XFILL_6_DFFSR_32 gnd vdd FILL
XFILL_6_DFFSR_43 gnd vdd FILL
XFILL_49_5_2 gnd vdd FILL
XFILL_69_DFFSR_114 gnd vdd FILL
XFILL_8_MUX2X1_38 gnd vdd FILL
XFILL_56_DFFSR_7 gnd vdd FILL
XFILL_8_MUX2X1_49 gnd vdd FILL
XFILL_6_DFFSR_54 gnd vdd FILL
XFILL_69_DFFSR_125 gnd vdd FILL
XFILL_32_DFFSR_40 gnd vdd FILL
XFILL_48_0_1 gnd vdd FILL
XFILL_6_DFFSR_65 gnd vdd FILL
XFILL_69_DFFSR_136 gnd vdd FILL
XFILL_6_DFFSR_76 gnd vdd FILL
XFILL_0_AOI22X1_1 gnd vdd FILL
XFILL_12_OAI21X1_4 gnd vdd FILL
XFILL_32_DFFSR_51 gnd vdd FILL
XFILL_69_DFFSR_147 gnd vdd FILL
XFILL_69_DFFSR_158 gnd vdd FILL
XFILL_6_DFFSR_87 gnd vdd FILL
XFILL_32_DFFSR_62 gnd vdd FILL
XFILL_6_DFFSR_98 gnd vdd FILL
XFILL_7_OAI22X1_30 gnd vdd FILL
XFILL_32_DFFSR_73 gnd vdd FILL
XFILL_69_DFFSR_169 gnd vdd FILL
XFILL_32_DFFSR_84 gnd vdd FILL
XFILL_7_OAI22X1_41 gnd vdd FILL
XFILL_32_DFFSR_95 gnd vdd FILL
XFILL_0_INVX1_200 gnd vdd FILL
XFILL_0_INVX1_211 gnd vdd FILL
XFILL_0_INVX1_222 gnd vdd FILL
XFILL_72_DFFSR_50 gnd vdd FILL
XFILL_72_DFFSR_61 gnd vdd FILL
XFILL_72_DFFSR_72 gnd vdd FILL
XFILL_72_DFFSR_83 gnd vdd FILL
XFILL_23_DFFSR_270 gnd vdd FILL
XFILL_72_DFFSR_94 gnd vdd FILL
XFILL_60_7_0 gnd vdd FILL
XFILL_20_MUX2X1_15 gnd vdd FILL
XFILL_4_INVX1_210 gnd vdd FILL
XFILL_32_4_2 gnd vdd FILL
XFILL_4_INVX1_221 gnd vdd FILL
XFILL_20_MUX2X1_26 gnd vdd FILL
XFILL_20_MUX2X1_37 gnd vdd FILL
XFILL_20_MUX2X1_48 gnd vdd FILL
XFILL_20_MUX2X1_59 gnd vdd FILL
XFILL_50_DFFSR_170 gnd vdd FILL
XFILL_12_NOR3X1_2 gnd vdd FILL
XFILL_0_OAI21X1_10 gnd vdd FILL
XFILL_0_OAI21X1_21 gnd vdd FILL
XFILL_41_DFFSR_60 gnd vdd FILL
XFILL_50_DFFSR_181 gnd vdd FILL
XFILL_50_DFFSR_192 gnd vdd FILL
XFILL_0_OAI21X1_32 gnd vdd FILL
XFILL_41_DFFSR_71 gnd vdd FILL
XFILL_41_DFFSR_82 gnd vdd FILL
XFILL_0_OAI21X1_43 gnd vdd FILL
XFILL_41_DFFSR_93 gnd vdd FILL
XFILL_54_DFFSR_180 gnd vdd FILL
XFILL_81_DFFSR_70 gnd vdd FILL
XFILL_54_DFFSR_191 gnd vdd FILL
XFILL_13_AOI21X1_80 gnd vdd FILL
XFILL_81_DFFSR_81 gnd vdd FILL
XFILL_81_DFFSR_92 gnd vdd FILL
XFILL_10_DFFSR_70 gnd vdd FILL
XFILL_10_DFFSR_81 gnd vdd FILL
XFILL_10_DFFSR_92 gnd vdd FILL
XFILL_32_DFFSR_104 gnd vdd FILL
XFILL_58_DFFSR_190 gnd vdd FILL
XFILL_32_DFFSR_115 gnd vdd FILL
XFILL_32_DFFSR_126 gnd vdd FILL
XFILL_32_DFFSR_137 gnd vdd FILL
XFILL_1_DFFSR_150 gnd vdd FILL
XFILL_1_DFFSR_161 gnd vdd FILL
XFILL_32_DFFSR_148 gnd vdd FILL
XFILL_50_DFFSR_80 gnd vdd FILL
XFILL_1_DFFSR_172 gnd vdd FILL
XFILL_32_DFFSR_159 gnd vdd FILL
XFILL_21_11 gnd vdd FILL
XFILL_1_DFFSR_183 gnd vdd FILL
XFILL_50_DFFSR_91 gnd vdd FILL
XFILL_39_0_1 gnd vdd FILL
XFILL_1_DFFSR_194 gnd vdd FILL
XFILL_36_DFFSR_103 gnd vdd FILL
XFILL_36_DFFSR_114 gnd vdd FILL
XFILL_36_DFFSR_125 gnd vdd FILL
XFILL_2_NAND3X1_19 gnd vdd FILL
XFILL_36_DFFSR_136 gnd vdd FILL
XFILL_5_DFFSR_160 gnd vdd FILL
XFILL_36_DFFSR_147 gnd vdd FILL
XFILL_36_DFFSR_158 gnd vdd FILL
XFILL_5_DFFSR_171 gnd vdd FILL
XFILL_36_DFFSR_169 gnd vdd FILL
XFILL_5_DFFSR_182 gnd vdd FILL
XFILL_5_DFFSR_193 gnd vdd FILL
XFILL_9_NAND3X1_130 gnd vdd FILL
XFILL_4_NOR3X1_1 gnd vdd FILL
XFILL_51_7_0 gnd vdd FILL
XFILL_16_MUX2X1_130 gnd vdd FILL
XFILL_9_DFFSR_170 gnd vdd FILL
XFILL_23_4_2 gnd vdd FILL
XFILL_16_MUX2X1_141 gnd vdd FILL
XFILL_9_DFFSR_181 gnd vdd FILL
XFILL_16_MUX2X1_152 gnd vdd FILL
XFILL_16_MUX2X1_163 gnd vdd FILL
XFILL_13_MUX2X1_90 gnd vdd FILL
XFILL_9_DFFSR_192 gnd vdd FILL
XFILL_16_MUX2X1_174 gnd vdd FILL
XFILL_1_NOR3X1_50 gnd vdd FILL
XFILL_16_MUX2X1_185 gnd vdd FILL
XFILL_82_DFFSR_204 gnd vdd FILL
XFILL_82_DFFSR_215 gnd vdd FILL
XFILL_82_DFFSR_226 gnd vdd FILL
XFILL_82_DFFSR_237 gnd vdd FILL
XFILL_3_DFFSR_2 gnd vdd FILL
XFILL_82_DFFSR_248 gnd vdd FILL
XFILL_82_DFFSR_259 gnd vdd FILL
XFILL_73_DFFSR_1 gnd vdd FILL
XFILL_2_DFFSR_80 gnd vdd FILL
XFILL_86_DFFSR_203 gnd vdd FILL
XFILL_2_DFFSR_91 gnd vdd FILL
XFILL_86_DFFSR_214 gnd vdd FILL
XFILL_86_DFFSR_225 gnd vdd FILL
XFILL_86_DFFSR_236 gnd vdd FILL
XFILL_86_DFFSR_247 gnd vdd FILL
XFILL_86_DFFSR_258 gnd vdd FILL
XFILL_21_DFFSR_180 gnd vdd FILL
XFILL_86_DFFSR_269 gnd vdd FILL
XFILL_2_INVX1_120 gnd vdd FILL
XFILL_21_DFFSR_191 gnd vdd FILL
XFILL_11_BUFX2_6 gnd vdd FILL
XFILL_2_INVX1_131 gnd vdd FILL
XFILL_2_INVX1_142 gnd vdd FILL
XFILL_2_INVX1_153 gnd vdd FILL
XFILL_2_INVX1_164 gnd vdd FILL
XFILL_2_INVX1_175 gnd vdd FILL
XFILL_2_INVX1_186 gnd vdd FILL
XFILL_2_INVX1_197 gnd vdd FILL
XFILL_25_DFFSR_190 gnd vdd FILL
XFILL_6_INVX1_130 gnd vdd FILL
XFILL_6_5_2 gnd vdd FILL
XFILL_6_INVX1_141 gnd vdd FILL
XFILL_6_INVX1_152 gnd vdd FILL
XFILL_38_DFFSR_4 gnd vdd FILL
XFILL_5_0_1 gnd vdd FILL
XFILL_6_INVX1_163 gnd vdd FILL
XFILL_6_INVX1_174 gnd vdd FILL
XFILL_6_INVX1_185 gnd vdd FILL
XFILL_6_MUX2X1_180 gnd vdd FILL
XFILL_6_INVX1_196 gnd vdd FILL
XFILL_6_MUX2X1_191 gnd vdd FILL
XFILL_0_OAI22X1_4 gnd vdd FILL
XFILL_42_7_0 gnd vdd FILL
XFILL_14_4_2 gnd vdd FILL
XFILL_2_NOR2X1_109 gnd vdd FILL
XFILL_4_OAI22X1_3 gnd vdd FILL
XFILL_8_OAI22X1_2 gnd vdd FILL
XFILL_53_DFFSR_203 gnd vdd FILL
XFILL_53_DFFSR_214 gnd vdd FILL
XFILL_53_DFFSR_225 gnd vdd FILL
XFILL_53_DFFSR_236 gnd vdd FILL
XFILL_9_NAND3X1_50 gnd vdd FILL
XFILL_53_DFFSR_247 gnd vdd FILL
XFILL_9_NAND3X1_61 gnd vdd FILL
XFILL_53_DFFSR_258 gnd vdd FILL
XFILL_53_DFFSR_269 gnd vdd FILL
XFILL_9_NAND3X1_72 gnd vdd FILL
XFILL_15_BUFX4_30 gnd vdd FILL
XFILL_80_DFFSR_103 gnd vdd FILL
XFILL_9_NAND3X1_83 gnd vdd FILL
XFILL_57_DFFSR_202 gnd vdd FILL
XFILL_9_NAND3X1_94 gnd vdd FILL
XFILL_15_BUFX4_41 gnd vdd FILL
XFILL_80_DFFSR_114 gnd vdd FILL
XFILL_57_DFFSR_213 gnd vdd FILL
XFILL_15_BUFX4_52 gnd vdd FILL
XFILL_1_4 gnd vdd FILL
XFILL_57_DFFSR_224 gnd vdd FILL
XFILL_80_DFFSR_125 gnd vdd FILL
XFILL_80_DFFSR_136 gnd vdd FILL
XFILL_57_DFFSR_235 gnd vdd FILL
XFILL_15_BUFX4_63 gnd vdd FILL
XFILL_15_BUFX4_74 gnd vdd FILL
XFILL_57_DFFSR_246 gnd vdd FILL
XFILL_80_DFFSR_147 gnd vdd FILL
XFILL_80_DFFSR_158 gnd vdd FILL
XFILL_15_BUFX4_85 gnd vdd FILL
XFILL_15_BUFX4_96 gnd vdd FILL
XFILL_80_DFFSR_169 gnd vdd FILL
XFILL_57_DFFSR_257 gnd vdd FILL
XFILL_57_DFFSR_268 gnd vdd FILL
XFILL_12_CLKBUF1_9 gnd vdd FILL
XFILL_0_DFFSR_206 gnd vdd FILL
XFILL_84_DFFSR_102 gnd vdd FILL
XFILL_12_AOI22X1_11 gnd vdd FILL
XFILL_64_DFFSR_19 gnd vdd FILL
XFILL_0_DFFSR_217 gnd vdd FILL
XFILL_84_DFFSR_113 gnd vdd FILL
XFILL_84_DFFSR_124 gnd vdd FILL
XFILL_0_DFFSR_228 gnd vdd FILL
XFILL_50_5 gnd vdd FILL
XFILL_84_DFFSR_135 gnd vdd FILL
XFILL_0_DFFSR_239 gnd vdd FILL
XFILL_84_DFFSR_146 gnd vdd FILL
XFILL_84_DFFSR_157 gnd vdd FILL
XFILL_64_3_2 gnd vdd FILL
XFILL_43_4 gnd vdd FILL
XFILL_84_DFFSR_168 gnd vdd FILL
XFILL_84_DFFSR_179 gnd vdd FILL
XFILL_2_NAND2X1_30 gnd vdd FILL
XFILL_16_CLKBUF1_8 gnd vdd FILL
XFILL_2_NAND2X1_41 gnd vdd FILL
XFILL_4_DFFSR_205 gnd vdd FILL
XFILL_1_NAND3X1_5 gnd vdd FILL
XFILL_2_NAND2X1_52 gnd vdd FILL
XFILL_4_DFFSR_216 gnd vdd FILL
XFILL_2_NAND2X1_63 gnd vdd FILL
XFILL_4_DFFSR_227 gnd vdd FILL
XFILL_2_NAND2X1_74 gnd vdd FILL
XFILL_4_DFFSR_238 gnd vdd FILL
XFILL_2_NAND2X1_85 gnd vdd FILL
XFILL_4_DFFSR_249 gnd vdd FILL
XFILL_2_NAND2X1_96 gnd vdd FILL
XFILL_33_7_0 gnd vdd FILL
XFILL_33_DFFSR_18 gnd vdd FILL
XFILL_12_BUFX4_103 gnd vdd FILL
XFILL_33_DFFSR_29 gnd vdd FILL
XFILL_10_CLKBUF1_16 gnd vdd FILL
XFILL_8_DFFSR_204 gnd vdd FILL
XFILL_5_NAND3X1_4 gnd vdd FILL
XFILL_8_DFFSR_215 gnd vdd FILL
XFILL_10_CLKBUF1_27 gnd vdd FILL
XFILL_8_DFFSR_226 gnd vdd FILL
XFILL_10_CLKBUF1_38 gnd vdd FILL
XFILL_8_DFFSR_237 gnd vdd FILL
XFILL_8_DFFSR_248 gnd vdd FILL
XFILL_73_DFFSR_17 gnd vdd FILL
XFILL_8_DFFSR_259 gnd vdd FILL
XFILL_73_DFFSR_28 gnd vdd FILL
XFILL_73_DFFSR_39 gnd vdd FILL
XFILL_9_NAND3X1_3 gnd vdd FILL
XFILL_16_MUX2X1_7 gnd vdd FILL
XFILL_16_11 gnd vdd FILL
XFILL_28_CLKBUF1_40 gnd vdd FILL
XFILL_7_BUFX4_40 gnd vdd FILL
XFILL_7_BUFX4_51 gnd vdd FILL
XFILL_7_BUFX4_62 gnd vdd FILL
XFILL_42_DFFSR_16 gnd vdd FILL
XFILL_7_BUFX4_73 gnd vdd FILL
XFILL_20_DFFSR_203 gnd vdd FILL
XFILL_42_DFFSR_27 gnd vdd FILL
XFILL_7_BUFX4_84 gnd vdd FILL
XFILL_42_DFFSR_38 gnd vdd FILL
XFILL_20_DFFSR_214 gnd vdd FILL
XFILL_19_MUX2X1_107 gnd vdd FILL
XFILL_10_NOR2X1_16 gnd vdd FILL
XFILL_7_BUFX4_95 gnd vdd FILL
XFILL_19_MUX2X1_118 gnd vdd FILL
XFILL_42_DFFSR_49 gnd vdd FILL
XFILL_20_DFFSR_225 gnd vdd FILL
XFILL_19_MUX2X1_129 gnd vdd FILL
XFILL_6_AOI21X1_30 gnd vdd FILL
XFILL_10_NOR2X1_27 gnd vdd FILL
XFILL_20_DFFSR_236 gnd vdd FILL
XFILL_6_AOI21X1_41 gnd vdd FILL
XFILL_32_10 gnd vdd FILL
XFILL_10_NOR2X1_38 gnd vdd FILL
XFILL_6_AOI21X1_52 gnd vdd FILL
XFILL_20_DFFSR_247 gnd vdd FILL
XFILL_10_NOR2X1_49 gnd vdd FILL
XFILL_20_DFFSR_258 gnd vdd FILL
XFILL_16_OAI22X1_10 gnd vdd FILL
XFILL_20_DFFSR_269 gnd vdd FILL
XFILL_6_AOI21X1_63 gnd vdd FILL
XFILL_16_OAI22X1_21 gnd vdd FILL
XFILL_6_AOI21X1_74 gnd vdd FILL
XFILL_16_OAI22X1_32 gnd vdd FILL
XFILL_1_INVX1_209 gnd vdd FILL
XFILL_82_DFFSR_15 gnd vdd FILL
XFILL_24_DFFSR_202 gnd vdd FILL
XFILL_16_OAI22X1_43 gnd vdd FILL
XFILL_82_DFFSR_26 gnd vdd FILL
XFILL_24_DFFSR_213 gnd vdd FILL
XFILL_82_DFFSR_37 gnd vdd FILL
XFILL_82_DFFSR_48 gnd vdd FILL
XFILL_24_DFFSR_224 gnd vdd FILL
XFILL_24_DFFSR_235 gnd vdd FILL
XFILL_5_AOI22X1_9 gnd vdd FILL
XFILL_82_DFFSR_59 gnd vdd FILL
XFILL_7_DFFSR_3 gnd vdd FILL
XFILL_9_NOR2X1_140 gnd vdd FILL
XFILL_11_DFFSR_15 gnd vdd FILL
XFILL_24_DFFSR_246 gnd vdd FILL
XFILL_11_DFFSR_26 gnd vdd FILL
XFILL_0_CLKBUF1_11 gnd vdd FILL
XFILL_11_DFFSR_37 gnd vdd FILL
XFILL_9_NOR2X1_151 gnd vdd FILL
XFILL_24_DFFSR_257 gnd vdd FILL
XFILL_0_CLKBUF1_22 gnd vdd FILL
XFILL_24_DFFSR_268 gnd vdd FILL
XFILL_9_NOR2X1_162 gnd vdd FILL
XFILL_11_DFFSR_48 gnd vdd FILL
XFILL_9_NOR2X1_173 gnd vdd FILL
XFILL_0_CLKBUF1_33 gnd vdd FILL
XFILL_77_DFFSR_2 gnd vdd FILL
XFILL_11_DFFSR_59 gnd vdd FILL
XFILL_28_DFFSR_201 gnd vdd FILL
XFILL_5_INVX1_208 gnd vdd FILL
XFILL_51_DFFSR_102 gnd vdd FILL
XFILL_9_NOR2X1_184 gnd vdd FILL
XFILL_55_3_2 gnd vdd FILL
XFILL_9_NOR2X1_8 gnd vdd FILL
XFILL_5_INVX1_219 gnd vdd FILL
XFILL_51_DFFSR_113 gnd vdd FILL
XFILL_51_DFFSR_124 gnd vdd FILL
XFILL_28_DFFSR_212 gnd vdd FILL
XFILL_9_NOR2X1_195 gnd vdd FILL
XFILL_28_DFFSR_223 gnd vdd FILL
XFILL_28_DFFSR_234 gnd vdd FILL
XFILL_51_DFFSR_135 gnd vdd FILL
XFILL_51_DFFSR_14 gnd vdd FILL
XFILL_9_AOI22X1_8 gnd vdd FILL
XFILL_51_DFFSR_146 gnd vdd FILL
XFILL_28_DFFSR_245 gnd vdd FILL
XFILL_51_DFFSR_157 gnd vdd FILL
XFILL_51_DFFSR_25 gnd vdd FILL
XFILL_51_DFFSR_36 gnd vdd FILL
XFILL_51_DFFSR_168 gnd vdd FILL
XFILL_28_DFFSR_256 gnd vdd FILL
XFILL_2_BUFX2_9 gnd vdd FILL
XFILL_28_DFFSR_267 gnd vdd FILL
XFILL_51_DFFSR_47 gnd vdd FILL
XFILL_51_DFFSR_179 gnd vdd FILL
XFILL_51_DFFSR_58 gnd vdd FILL
XFILL_55_DFFSR_101 gnd vdd FILL
XFILL_51_DFFSR_69 gnd vdd FILL
XFILL_24_7_0 gnd vdd FILL
XFILL_55_DFFSR_112 gnd vdd FILL
XFILL_55_DFFSR_123 gnd vdd FILL
XFILL_55_DFFSR_134 gnd vdd FILL
XFILL_55_DFFSR_145 gnd vdd FILL
XFILL_55_DFFSR_156 gnd vdd FILL
XFILL_8_MUX2X1_6 gnd vdd FILL
XFILL_55_DFFSR_167 gnd vdd FILL
XFILL_55_DFFSR_178 gnd vdd FILL
XFILL_20_DFFSR_13 gnd vdd FILL
XFILL_9_MUX2X1_102 gnd vdd FILL
XFILL_20_DFFSR_24 gnd vdd FILL
XFILL_59_DFFSR_100 gnd vdd FILL
XFILL_55_DFFSR_189 gnd vdd FILL
XFILL_9_MUX2X1_113 gnd vdd FILL
XFILL_61_DFFSR_8 gnd vdd FILL
XFILL_59_DFFSR_111 gnd vdd FILL
XFILL_20_DFFSR_35 gnd vdd FILL
XFILL_9_MUX2X1_124 gnd vdd FILL
XFILL_59_DFFSR_122 gnd vdd FILL
XFILL_59_DFFSR_133 gnd vdd FILL
XFILL_20_DFFSR_46 gnd vdd FILL
XFILL_9_MUX2X1_135 gnd vdd FILL
XFILL_9_MUX2X1_146 gnd vdd FILL
XFILL_20_DFFSR_57 gnd vdd FILL
XFILL_59_DFFSR_144 gnd vdd FILL
XFILL_20_DFFSR_68 gnd vdd FILL
XFILL_59_DFFSR_155 gnd vdd FILL
XFILL_20_DFFSR_79 gnd vdd FILL
XFILL_9_MUX2X1_157 gnd vdd FILL
XFILL_9_MUX2X1_168 gnd vdd FILL
XFILL_59_DFFSR_166 gnd vdd FILL
XFILL_59_DFFSR_177 gnd vdd FILL
XFILL_9_MUX2X1_179 gnd vdd FILL
XFILL_2_DFFSR_104 gnd vdd FILL
XFILL_60_DFFSR_12 gnd vdd FILL
XFILL_59_DFFSR_188 gnd vdd FILL
XFILL_2_DFFSR_115 gnd vdd FILL
XFILL_60_DFFSR_23 gnd vdd FILL
XFILL_60_DFFSR_34 gnd vdd FILL
XFILL_59_DFFSR_199 gnd vdd FILL
XFILL_31_NOR3X1_9 gnd vdd FILL
XFILL_2_DFFSR_126 gnd vdd FILL
XFILL_2_DFFSR_137 gnd vdd FILL
XFILL_60_DFFSR_45 gnd vdd FILL
XFILL_60_DFFSR_56 gnd vdd FILL
XFILL_2_DFFSR_148 gnd vdd FILL
XFILL_60_DFFSR_67 gnd vdd FILL
XDFFSR_70 DFFSR_70/Q DFFSR_70/CLK DFFSR_84/R vdd DFFSR_70/D gnd vdd DFFSR
XFILL_2_DFFSR_159 gnd vdd FILL
XFILL_60_DFFSR_78 gnd vdd FILL
XDFFSR_81 DFFSR_81/Q DFFSR_81/CLK DFFSR_84/R vdd DFFSR_81/D gnd vdd DFFSR
XFILL_60_DFFSR_89 gnd vdd FILL
XDFFSR_92 DFFSR_92/Q DFFSR_93/CLK DFFSR_93/R vdd DFFSR_92/D gnd vdd DFFSR
XFILL_6_DFFSR_103 gnd vdd FILL
XFILL_6_DFFSR_114 gnd vdd FILL
XFILL_10_MUX2X1_12 gnd vdd FILL
XFILL_10_MUX2X1_23 gnd vdd FILL
XFILL_3_DFFSR_14 gnd vdd FILL
XFILL_6_DFFSR_125 gnd vdd FILL
XFILL_3_DFFSR_25 gnd vdd FILL
XFILL_6_DFFSR_136 gnd vdd FILL
XFILL_1_BUFX4_3 gnd vdd FILL
XFILL_10_MUX2X1_34 gnd vdd FILL
XFILL_3_DFFSR_36 gnd vdd FILL
XFILL_10_MUX2X1_45 gnd vdd FILL
XFILL_6_DFFSR_147 gnd vdd FILL
XFILL_6_DFFSR_158 gnd vdd FILL
XFILL_10_MUX2X1_56 gnd vdd FILL
XFILL_3_DFFSR_47 gnd vdd FILL
XFILL_3_DFFSR_58 gnd vdd FILL
XFILL_14_BUFX4_1 gnd vdd FILL
XFILL_6_DFFSR_169 gnd vdd FILL
XFILL_10_MUX2X1_67 gnd vdd FILL
XFILL_10_MUX2X1_78 gnd vdd FILL
XFILL_3_DFFSR_69 gnd vdd FILL
XFILL_10_MUX2X1_89 gnd vdd FILL
XFILL_14_MUX2X1_11 gnd vdd FILL
XFILL_14_MUX2X1_22 gnd vdd FILL
XFILL_14_MUX2X1_33 gnd vdd FILL
XFILL_5_INVX1_90 gnd vdd FILL
XFILL_14_MUX2X1_44 gnd vdd FILL
XFILL_5_BUFX2_10 gnd vdd FILL
XFILL_14_MUX2X1_55 gnd vdd FILL
XFILL_14_MUX2X1_66 gnd vdd FILL
XFILL_14_MUX2X1_77 gnd vdd FILL
XFILL_46_3_2 gnd vdd FILL
XFILL_2_NOR3X1_15 gnd vdd FILL
XFILL_14_MUX2X1_88 gnd vdd FILL
XFILL_2_NOR3X1_26 gnd vdd FILL
XFILL_14_MUX2X1_99 gnd vdd FILL
XFILL_18_MUX2X1_10 gnd vdd FILL
XFILL_2_NOR3X1_37 gnd vdd FILL
XFILL_18_MUX2X1_21 gnd vdd FILL
XFILL_2_NOR3X1_48 gnd vdd FILL
XFILL_18_MUX2X1_32 gnd vdd FILL
XFILL_18_MUX2X1_43 gnd vdd FILL
XFILL_18_MUX2X1_54 gnd vdd FILL
XFILL_18_MUX2X1_65 gnd vdd FILL
XFILL_15_7_0 gnd vdd FILL
XFILL_0_INVX1_7 gnd vdd FILL
XFILL_18_MUX2X1_76 gnd vdd FILL
XFILL_18_MUX2X1_87 gnd vdd FILL
XFILL_6_NOR3X1_14 gnd vdd FILL
XFILL_22_9 gnd vdd FILL
XFILL_6_NOR3X1_25 gnd vdd FILL
XFILL_6_NOR3X1_36 gnd vdd FILL
XFILL_18_MUX2X1_98 gnd vdd FILL
XFILL_22_DFFSR_101 gnd vdd FILL
XFILL_6_NOR3X1_47 gnd vdd FILL
XFILL_22_DFFSR_112 gnd vdd FILL
XFILL_22_DFFSR_123 gnd vdd FILL
XFILL_22_DFFSR_134 gnd vdd FILL
XFILL_22_DFFSR_145 gnd vdd FILL
XFILL_22_DFFSR_156 gnd vdd FILL
XFILL_22_DFFSR_167 gnd vdd FILL
XFILL_22_DFFSR_178 gnd vdd FILL
XFILL_3_INVX1_107 gnd vdd FILL
XFILL_3_INVX1_118 gnd vdd FILL
XFILL_26_DFFSR_100 gnd vdd FILL
XFILL_22_DFFSR_189 gnd vdd FILL
XFILL_26_DFFSR_111 gnd vdd FILL
XFILL_3_INVX1_129 gnd vdd FILL
XFILL_1_NAND3X1_16 gnd vdd FILL
XFILL_26_DFFSR_122 gnd vdd FILL
XFILL_26_DFFSR_133 gnd vdd FILL
XFILL_1_NAND3X1_27 gnd vdd FILL
XFILL_26_DFFSR_144 gnd vdd FILL
XFILL_1_NAND3X1_38 gnd vdd FILL
XFILL_26_DFFSR_155 gnd vdd FILL
XFILL_1_NAND3X1_49 gnd vdd FILL
XFILL_26_DFFSR_166 gnd vdd FILL
XFILL_26_DFFSR_177 gnd vdd FILL
XFILL_5_NAND2X1_18 gnd vdd FILL
XFILL_7_INVX1_106 gnd vdd FILL
XINVX1_120 INVX1_120/A gnd INVX1_120/Y vdd INVX1
XFILL_5_NAND2X1_29 gnd vdd FILL
XFILL_5_NOR2X1_1 gnd vdd FILL
XFILL_7_INVX1_117 gnd vdd FILL
XFILL_26_DFFSR_188 gnd vdd FILL
XINVX1_131 INVX1_131/A gnd INVX1_131/Y vdd INVX1
XFILL_7_INVX1_128 gnd vdd FILL
XFILL_26_DFFSR_199 gnd vdd FILL
XINVX1_142 BUFX2_7/A gnd NOR2X1_13/B vdd INVX1
XINVX1_153 INVX1_153/A gnd INVX1_153/Y vdd INVX1
XFILL_4_INVX8_1 gnd vdd FILL
XFILL_7_INVX1_139 gnd vdd FILL
XINVX1_164 INVX1_164/A gnd INVX1_164/Y vdd INVX1
XINVX1_175 INVX1_175/A gnd INVX1_175/Y vdd INVX1
XINVX1_186 INVX1_186/A gnd INVX1_186/Y vdd INVX1
XINVX1_197 DFFSR_89/Q gnd INVX1_197/Y vdd INVX1
XFILL_29_DFFSR_90 gnd vdd FILL
XFILL_22_NOR3X1_12 gnd vdd FILL
XFILL_15_MUX2X1_160 gnd vdd FILL
XFILL_15_MUX2X1_171 gnd vdd FILL
XFILL_22_NOR3X1_23 gnd vdd FILL
XFILL_22_NOR3X1_34 gnd vdd FILL
XFILL_15_MUX2X1_182 gnd vdd FILL
XFILL_22_NOR3X1_45 gnd vdd FILL
XFILL_72_DFFSR_201 gnd vdd FILL
XFILL_15_MUX2X1_193 gnd vdd FILL
XFILL_72_DFFSR_212 gnd vdd FILL
XFILL_72_DFFSR_223 gnd vdd FILL
XFILL_72_DFFSR_234 gnd vdd FILL
XFILL_72_DFFSR_245 gnd vdd FILL
XFILL_26_NOR3X1_11 gnd vdd FILL
XFILL_21_DFFSR_1 gnd vdd FILL
XFILL_72_DFFSR_256 gnd vdd FILL
XFILL_72_DFFSR_267 gnd vdd FILL
XFILL_26_NOR3X1_22 gnd vdd FILL
XFILL_26_NOR3X1_33 gnd vdd FILL
XFILL_65_6_0 gnd vdd FILL
XFILL_76_DFFSR_200 gnd vdd FILL
XFILL_26_NOR3X1_44 gnd vdd FILL
XFILL_37_3_2 gnd vdd FILL
XFILL_76_DFFSR_211 gnd vdd FILL
XFILL_76_DFFSR_222 gnd vdd FILL
XFILL_76_DFFSR_233 gnd vdd FILL
XFILL_76_DFFSR_244 gnd vdd FILL
XFILL_1_NOR3X1_5 gnd vdd FILL
XFILL_76_DFFSR_255 gnd vdd FILL
XFILL_76_DFFSR_266 gnd vdd FILL
XFILL_31_CLKBUF1_7 gnd vdd FILL
XFILL_9_AOI21X1_18 gnd vdd FILL
XFILL_9_AOI21X1_29 gnd vdd FILL
XFILL_35_CLKBUF1_6 gnd vdd FILL
XFILL_20_CLKBUF1_17 gnd vdd FILL
XFILL_20_CLKBUF1_28 gnd vdd FILL
XFILL_20_2_2 gnd vdd FILL
XFILL_27_10 gnd vdd FILL
XFILL_43_DFFSR_5 gnd vdd FILL
XFILL_20_CLKBUF1_39 gnd vdd FILL
XFILL_1_NOR2X1_106 gnd vdd FILL
XFILL_1_NOR2X1_117 gnd vdd FILL
XFILL_1_NOR2X1_128 gnd vdd FILL
XFILL_1_NOR2X1_139 gnd vdd FILL
XFILL_11_NAND2X1_10 gnd vdd FILL
XFILL_65_DFFSR_9 gnd vdd FILL
XFILL_11_NAND2X1_21 gnd vdd FILL
XFILL_8_BUFX4_18 gnd vdd FILL
XFILL_11_NAND2X1_32 gnd vdd FILL
XFILL_8_BUFX4_29 gnd vdd FILL
XFILL_11_NAND2X1_43 gnd vdd FILL
XFILL_1_OAI21X1_2 gnd vdd FILL
XFILL_11_NAND2X1_54 gnd vdd FILL
XFILL_11_NAND2X1_65 gnd vdd FILL
XFILL_56_6_0 gnd vdd FILL
XFILL_9_OAI22X1_15 gnd vdd FILL
XFILL_11_NAND2X1_76 gnd vdd FILL
XFILL_9_OAI22X1_26 gnd vdd FILL
XFILL_28_3_2 gnd vdd FILL
XFILL_3_3_2 gnd vdd FILL
XFILL_11_NAND2X1_87 gnd vdd FILL
XFILL_9_OAI22X1_37 gnd vdd FILL
XFILL_9_OAI22X1_48 gnd vdd FILL
XFILL_43_DFFSR_200 gnd vdd FILL
XFILL_43_DFFSR_211 gnd vdd FILL
XFILL_43_DFFSR_222 gnd vdd FILL
XFILL_5_OAI21X1_1 gnd vdd FILL
XFILL_43_DFFSR_233 gnd vdd FILL
XFILL_43_DFFSR_244 gnd vdd FILL
XFILL_43_DFFSR_255 gnd vdd FILL
XFILL_2_NOR2X1_70 gnd vdd FILL
XFILL_2_NOR2X1_81 gnd vdd FILL
XFILL_43_DFFSR_266 gnd vdd FILL
XNAND3X1_106 NAND3X1_106/A NAND3X1_106/B NAND3X1_106/C gnd NOR3X1_28/C vdd NAND3X1
XFILL_2_NOR2X1_92 gnd vdd FILL
XNAND3X1_117 NOR2X1_2/A BUFX4_91/Y NOR2X1_37/Y gnd NAND3X1_118/C vdd NAND3X1
XFILL_8_NAND3X1_80 gnd vdd FILL
XNAND3X1_128 INVX1_162/A BUFX4_90/Y NOR3X1_51/Y gnd OAI21X1_20/C vdd NAND3X1
XFILL_70_DFFSR_100 gnd vdd FILL
XFILL_8_NAND3X1_91 gnd vdd FILL
XFILL_70_DFFSR_111 gnd vdd FILL
XFILL_5_BUFX4_4 gnd vdd FILL
XFILL_47_DFFSR_210 gnd vdd FILL
XFILL_70_DFFSR_122 gnd vdd FILL
XFILL_6_NOR2X1_206 gnd vdd FILL
XFILL_47_DFFSR_221 gnd vdd FILL
XFILL_70_DFFSR_133 gnd vdd FILL
XFILL_47_DFFSR_232 gnd vdd FILL
XFILL_47_DFFSR_243 gnd vdd FILL
XFILL_70_DFFSR_144 gnd vdd FILL
XFILL_70_DFFSR_155 gnd vdd FILL
XFILL_47_DFFSR_254 gnd vdd FILL
XFILL_11_2_2 gnd vdd FILL
XFILL_70_DFFSR_166 gnd vdd FILL
XFILL_70_DFFSR_177 gnd vdd FILL
XFILL_6_NOR2X1_80 gnd vdd FILL
XFILL_47_DFFSR_265 gnd vdd FILL
XFILL_15_AND2X2_6 gnd vdd FILL
XFILL_2_OAI21X1_17 gnd vdd FILL
XFILL_6_NOR2X1_91 gnd vdd FILL
XFILL_2_OAI21X1_28 gnd vdd FILL
XFILL_70_DFFSR_188 gnd vdd FILL
XFILL_74_DFFSR_110 gnd vdd FILL
XFILL_70_DFFSR_199 gnd vdd FILL
XFILL_74_DFFSR_121 gnd vdd FILL
XFILL_2_OAI21X1_39 gnd vdd FILL
XFILL_74_DFFSR_132 gnd vdd FILL
XFILL_74_DFFSR_143 gnd vdd FILL
XFILL_15_AOI21X1_10 gnd vdd FILL
XFILL_74_DFFSR_154 gnd vdd FILL
XFILL_15_AOI21X1_21 gnd vdd FILL
XFILL_15_AOI21X1_32 gnd vdd FILL
XFILL_74_DFFSR_165 gnd vdd FILL
XFILL_74_DFFSR_176 gnd vdd FILL
XFILL_15_AOI21X1_43 gnd vdd FILL
XFILL_74_DFFSR_187 gnd vdd FILL
XFILL_15_AOI21X1_54 gnd vdd FILL
XFILL_74_DFFSR_198 gnd vdd FILL
XFILL_15_AOI21X1_65 gnd vdd FILL
XFILL_12_BUFX4_12 gnd vdd FILL
XFILL_1_NAND2X1_60 gnd vdd FILL
XFILL_78_DFFSR_120 gnd vdd FILL
XFILL_15_AOI21X1_76 gnd vdd FILL
XFILL_78_DFFSR_131 gnd vdd FILL
XFILL_12_BUFX4_23 gnd vdd FILL
XFILL_1_NAND2X1_71 gnd vdd FILL
XFILL_78_DFFSR_142 gnd vdd FILL
XFILL_1_NAND2X1_82 gnd vdd FILL
XFILL_12_BUFX4_34 gnd vdd FILL
XFILL_4_INVX1_8 gnd vdd FILL
XFILL_12_BUFX4_45 gnd vdd FILL
XFILL_1_NAND2X1_93 gnd vdd FILL
XFILL_78_DFFSR_153 gnd vdd FILL
XFILL_12_BUFX4_56 gnd vdd FILL
XFILL_78_DFFSR_164 gnd vdd FILL
XFILL_78_DFFSR_175 gnd vdd FILL
XFILL_12_BUFX4_67 gnd vdd FILL
XFILL_12_BUFX4_78 gnd vdd FILL
XFILL_78_DFFSR_186 gnd vdd FILL
XFILL_12_BUFX4_89 gnd vdd FILL
XFILL_78_DFFSR_197 gnd vdd FILL
XFILL_2_NAND2X1_3 gnd vdd FILL
XFILL_47_6_0 gnd vdd FILL
XFILL_19_3_2 gnd vdd FILL
XFILL_6_INVX1_13 gnd vdd FILL
XFILL_6_NAND2X1_2 gnd vdd FILL
XFILL_6_INVX1_24 gnd vdd FILL
XFILL_10_DFFSR_200 gnd vdd FILL
XFILL_61_1_2 gnd vdd FILL
XFILL_10_DFFSR_211 gnd vdd FILL
XFILL_6_INVX1_35 gnd vdd FILL
XFILL_8_INVX8_2 gnd vdd FILL
XFILL_18_MUX2X1_104 gnd vdd FILL
XFILL_6_INVX1_46 gnd vdd FILL
XFILL_10_DFFSR_222 gnd vdd FILL
XFILL_18_MUX2X1_115 gnd vdd FILL
XFILL_7_AND2X2_5 gnd vdd FILL
XFILL_10_DFFSR_233 gnd vdd FILL
XFILL_18_MUX2X1_126 gnd vdd FILL
XFILL_6_INVX1_57 gnd vdd FILL
XFILL_18_MUX2X1_137 gnd vdd FILL
XFILL_10_DFFSR_244 gnd vdd FILL
XFILL_6_INVX1_68 gnd vdd FILL
XFILL_10_DFFSR_255 gnd vdd FILL
XFILL_18_MUX2X1_148 gnd vdd FILL
XFILL_6_INVX1_79 gnd vdd FILL
XFILL_18_MUX2X1_159 gnd vdd FILL
XFILL_5_AOI21X1_60 gnd vdd FILL
XFILL_10_DFFSR_266 gnd vdd FILL
XFILL_5_AOI21X1_71 gnd vdd FILL
XFILL_13_5 gnd vdd FILL
XFILL_15_OAI22X1_40 gnd vdd FILL
XFILL_30_5_0 gnd vdd FILL
XFILL_15_OAI22X1_51 gnd vdd FILL
XFILL_14_DFFSR_210 gnd vdd FILL
XFILL_14_DFFSR_221 gnd vdd FILL
XFILL_14_DFFSR_232 gnd vdd FILL
XFILL_14_DFFSR_243 gnd vdd FILL
XFILL_25_DFFSR_2 gnd vdd FILL
XDFFSR_104 DFFSR_104/Q DFFSR_97/CLK DFFSR_97/R vdd DFFSR_104/D gnd vdd DFFSR
XFILL_4_BUFX4_11 gnd vdd FILL
XFILL_14_DFFSR_254 gnd vdd FILL
XDFFSR_115 INVX1_186/A DFFSR_52/CLK DFFSR_56/R vdd DFFSR_115/D gnd vdd DFFSR
XFILL_14_DFFSR_265 gnd vdd FILL
XFILL_82_DFFSR_3 gnd vdd FILL
XFILL_4_BUFX4_22 gnd vdd FILL
XDFFSR_126 INVX1_170/A DFFSR_2/CLK DFFSR_2/R vdd DFFSR_126/D gnd vdd DFFSR
XFILL_8_NOR2X1_170 gnd vdd FILL
XDFFSR_137 INVX1_162/A CLKBUF1_8/Y DFFSR_55/R vdd DFFSR_137/D gnd vdd DFFSR
XFILL_4_BUFX4_33 gnd vdd FILL
XFILL_8_NOR2X1_181 gnd vdd FILL
XDFFSR_148 DFFSR_148/Q CLKBUF1_6/Y DFFSR_48/R vdd DFFSR_148/D gnd vdd DFFSR
XFILL_4_BUFX4_44 gnd vdd FILL
XFILL_41_DFFSR_110 gnd vdd FILL
XFILL_8_NOR2X1_192 gnd vdd FILL
XFILL_41_DFFSR_121 gnd vdd FILL
XFILL_4_BUFX4_55 gnd vdd FILL
XFILL_18_DFFSR_220 gnd vdd FILL
XDFFSR_159 DFFSR_159/Q DFFSR_70/CLK DFFSR_96/R vdd DFFSR_159/D gnd vdd DFFSR
XFILL_4_BUFX4_66 gnd vdd FILL
XFILL_41_DFFSR_132 gnd vdd FILL
XFILL_2_AOI21X1_8 gnd vdd FILL
XFILL_18_DFFSR_231 gnd vdd FILL
XFILL_41_DFFSR_143 gnd vdd FILL
XFILL_18_DFFSR_242 gnd vdd FILL
XFILL_4_BUFX4_77 gnd vdd FILL
XFILL_41_DFFSR_154 gnd vdd FILL
XFILL_18_DFFSR_253 gnd vdd FILL
XFILL_4_BUFX4_88 gnd vdd FILL
XFILL_4_BUFX4_99 gnd vdd FILL
XFILL_41_DFFSR_165 gnd vdd FILL
XFILL_18_DFFSR_264 gnd vdd FILL
XFILL_41_DFFSR_176 gnd vdd FILL
XFILL_18_DFFSR_275 gnd vdd FILL
XFILL_41_DFFSR_187 gnd vdd FILL
XFILL_41_DFFSR_198 gnd vdd FILL
XFILL_45_DFFSR_120 gnd vdd FILL
XFILL_45_DFFSR_131 gnd vdd FILL
XFILL_6_AOI21X1_7 gnd vdd FILL
XFILL_45_DFFSR_142 gnd vdd FILL
XFILL_45_DFFSR_153 gnd vdd FILL
XFILL_45_DFFSR_164 gnd vdd FILL
XFILL_45_DFFSR_175 gnd vdd FILL
XFILL_22_MUX2X1_9 gnd vdd FILL
XFILL_45_DFFSR_186 gnd vdd FILL
XFILL_8_MUX2X1_110 gnd vdd FILL
XFILL_19_MUX2X1_19 gnd vdd FILL
XFILL_45_DFFSR_197 gnd vdd FILL
XFILL_8_MUX2X1_121 gnd vdd FILL
XFILL_49_DFFSR_130 gnd vdd FILL
XFILL_47_DFFSR_6 gnd vdd FILL
XFILL_8_MUX2X1_132 gnd vdd FILL
XFILL_8_MUX2X1_143 gnd vdd FILL
XFILL_49_DFFSR_141 gnd vdd FILL
XNOR3X1_15 NOR3X1_15/A NOR3X1_49/B NOR3X1_1/B gnd NOR3X1_17/A vdd NOR3X1
XFILL_8_MUX2X1_154 gnd vdd FILL
XFILL_49_DFFSR_152 gnd vdd FILL
XNOR3X1_26 NOR3X1_26/A NOR3X1_46/B NOR3X1_46/C gnd NOR3X1_27/A vdd NOR3X1
XFILL_38_6_0 gnd vdd FILL
XFILL_11_AOI22X1_4 gnd vdd FILL
XFILL_8_MUX2X1_165 gnd vdd FILL
XFILL_49_DFFSR_163 gnd vdd FILL
XFILL_49_DFFSR_174 gnd vdd FILL
XFILL_8_MUX2X1_176 gnd vdd FILL
XNOR3X1_37 INVX1_71/Y NOR3X1_1/B INVX2_2/Y gnd NOR3X1_38/A vdd NOR3X1
XFILL_8_MUX2X1_187 gnd vdd FILL
XNOR3X1_48 INVX2_3/Y NOR3X1_48/B NOR3X1_48/C gnd NOR3X1_48/Y vdd NOR3X1
XFILL_49_DFFSR_185 gnd vdd FILL
XFILL_49_DFFSR_196 gnd vdd FILL
XFILL_15_AOI22X1_3 gnd vdd FILL
XFILL_52_1_2 gnd vdd FILL
XFILL_27_DFFSR_109 gnd vdd FILL
XFILL_19_AOI22X1_2 gnd vdd FILL
XFILL_10_NAND3X1_18 gnd vdd FILL
XFILL_10_NAND3X1_29 gnd vdd FILL
XFILL_21_5_0 gnd vdd FILL
XFILL_39_DFFSR_11 gnd vdd FILL
XFILL_30_CLKBUF1_18 gnd vdd FILL
XFILL_39_DFFSR_22 gnd vdd FILL
XFILL_30_CLKBUF1_29 gnd vdd FILL
XFILL_39_DFFSR_33 gnd vdd FILL
XFILL_39_DFFSR_44 gnd vdd FILL
XFILL_39_DFFSR_55 gnd vdd FILL
XFILL_39_DFFSR_66 gnd vdd FILL
XFILL_39_DFFSR_77 gnd vdd FILL
XFILL_39_DFFSR_88 gnd vdd FILL
XFILL_39_DFFSR_99 gnd vdd FILL
XFILL_79_DFFSR_10 gnd vdd FILL
XFILL_79_DFFSR_21 gnd vdd FILL
XFILL_79_DFFSR_32 gnd vdd FILL
XFILL_79_DFFSR_43 gnd vdd FILL
XFILL_0_DFFSR_18 gnd vdd FILL
XFILL_79_DFFSR_54 gnd vdd FILL
XFILL_0_DFFSR_29 gnd vdd FILL
XFILL_10_NOR2X1_6 gnd vdd FILL
XFILL_79_DFFSR_65 gnd vdd FILL
XFILL_79_DFFSR_76 gnd vdd FILL
XFILL_79_DFFSR_87 gnd vdd FILL
XFILL_79_DFFSR_98 gnd vdd FILL
XFILL_12_DFFSR_120 gnd vdd FILL
XFILL_2_INVX1_50 gnd vdd FILL
XFILL_9_BUFX4_5 gnd vdd FILL
XFILL_12_DFFSR_131 gnd vdd FILL
XFILL_2_INVX1_61 gnd vdd FILL
XFILL_77_DFFSR_209 gnd vdd FILL
XFILL_2_INVX1_72 gnd vdd FILL
XFILL_12_DFFSR_142 gnd vdd FILL
XFILL_2_INVX1_83 gnd vdd FILL
XFILL_2_INVX1_94 gnd vdd FILL
XFILL_12_DFFSR_153 gnd vdd FILL
XFILL_48_DFFSR_20 gnd vdd FILL
XFILL_48_DFFSR_31 gnd vdd FILL
XFILL_12_DFFSR_164 gnd vdd FILL
XFILL_12_DFFSR_175 gnd vdd FILL
XFILL_19_NOR3X1_6 gnd vdd FILL
XFILL_48_DFFSR_42 gnd vdd FILL
XFILL_1_CLKBUF1_7 gnd vdd FILL
XFILL_48_DFFSR_53 gnd vdd FILL
XFILL_12_DFFSR_186 gnd vdd FILL
XFILL_48_DFFSR_64 gnd vdd FILL
XFILL_12_DFFSR_197 gnd vdd FILL
XFILL_48_DFFSR_75 gnd vdd FILL
XFILL_0_NAND3X1_13 gnd vdd FILL
XFILL_29_6_0 gnd vdd FILL
XFILL_16_DFFSR_130 gnd vdd FILL
XFILL_48_DFFSR_86 gnd vdd FILL
XFILL_4_6_0 gnd vdd FILL
XFILL_0_NAND3X1_24 gnd vdd FILL
XFILL_16_DFFSR_141 gnd vdd FILL
XFILL_48_DFFSR_97 gnd vdd FILL
XFILL_0_NAND3X1_35 gnd vdd FILL
XFILL_16_DFFSR_152 gnd vdd FILL
XFILL_0_NAND3X1_46 gnd vdd FILL
XFILL_0_NAND3X1_57 gnd vdd FILL
XFILL_16_DFFSR_163 gnd vdd FILL
XFILL_16_DFFSR_174 gnd vdd FILL
XFILL_0_NAND3X1_68 gnd vdd FILL
XFILL_4_NAND2X1_15 gnd vdd FILL
XFILL_5_CLKBUF1_6 gnd vdd FILL
XFILL_4_NAND2X1_26 gnd vdd FILL
XFILL_16_DFFSR_185 gnd vdd FILL
XFILL_0_NAND3X1_79 gnd vdd FILL
XFILL_4_NAND2X1_37 gnd vdd FILL
XFILL_4_NAND2X1_48 gnd vdd FILL
XFILL_16_DFFSR_196 gnd vdd FILL
XFILL_0_BUFX4_70 gnd vdd FILL
XFILL_17_DFFSR_30 gnd vdd FILL
XFILL_0_BUFX4_81 gnd vdd FILL
XFILL_43_1_2 gnd vdd FILL
XFILL_4_NAND2X1_59 gnd vdd FILL
XFILL_17_DFFSR_41 gnd vdd FILL
XFILL_17_DFFSR_52 gnd vdd FILL
XFILL_17_DFFSR_63 gnd vdd FILL
XFILL_0_BUFX4_92 gnd vdd FILL
XFILL_1_BUFX4_101 gnd vdd FILL
XFILL_17_DFFSR_74 gnd vdd FILL
XFILL_17_DFFSR_85 gnd vdd FILL
XFILL_9_CLKBUF1_5 gnd vdd FILL
XFILL_17_DFFSR_96 gnd vdd FILL
XFILL_5_BUFX2_1 gnd vdd FILL
XFILL_12_NOR3X1_20 gnd vdd FILL
XFILL_12_NOR3X1_31 gnd vdd FILL
XFILL_14_MUX2X1_190 gnd vdd FILL
XFILL_12_5_0 gnd vdd FILL
XFILL_12_NOR3X1_42 gnd vdd FILL
XFILL_28_NOR3X1_4 gnd vdd FILL
XFILL_57_DFFSR_40 gnd vdd FILL
XFILL_57_DFFSR_51 gnd vdd FILL
XFILL_57_DFFSR_62 gnd vdd FILL
XFILL_62_DFFSR_220 gnd vdd FILL
XFILL_57_DFFSR_73 gnd vdd FILL
XFILL_62_DFFSR_231 gnd vdd FILL
XFILL_5_BUFX4_100 gnd vdd FILL
XFILL_57_DFFSR_84 gnd vdd FILL
XFILL_62_DFFSR_242 gnd vdd FILL
XFILL_62_DFFSR_253 gnd vdd FILL
XFILL_57_DFFSR_95 gnd vdd FILL
XFILL_62_DFFSR_264 gnd vdd FILL
XFILL_62_DFFSR_275 gnd vdd FILL
XFILL_16_NOR3X1_30 gnd vdd FILL
XFILL_16_NOR3X1_41 gnd vdd FILL
XFILL_16_NOR3X1_52 gnd vdd FILL
XFILL_2_NOR2X1_5 gnd vdd FILL
XFILL_10_NOR2X1_108 gnd vdd FILL
XFILL_66_DFFSR_230 gnd vdd FILL
XFILL_10_NOR2X1_119 gnd vdd FILL
XFILL_66_DFFSR_241 gnd vdd FILL
XFILL_66_DFFSR_252 gnd vdd FILL
XFILL_66_DFFSR_263 gnd vdd FILL
XFILL_26_DFFSR_50 gnd vdd FILL
XFILL_21_CLKBUF1_4 gnd vdd FILL
XFILL_26_DFFSR_61 gnd vdd FILL
XFILL_66_DFFSR_274 gnd vdd FILL
XFILL_26_DFFSR_72 gnd vdd FILL
XFILL_26_DFFSR_83 gnd vdd FILL
XFILL_26_DFFSR_94 gnd vdd FILL
XFILL_8_AOI21X1_15 gnd vdd FILL
XFILL_8_AOI21X1_26 gnd vdd FILL
XFILL_8_AOI21X1_37 gnd vdd FILL
XFILL_1_MUX2X1_3 gnd vdd FILL
XFILL_8_AOI21X1_48 gnd vdd FILL
XFILL_8_AOI21X1_59 gnd vdd FILL
XFILL_25_CLKBUF1_3 gnd vdd FILL
XFILL_18_OAI22X1_17 gnd vdd FILL
XFILL_66_DFFSR_60 gnd vdd FILL
XFILL_18_OAI22X1_28 gnd vdd FILL
XFILL_66_DFFSR_71 gnd vdd FILL
XFILL_66_DFFSR_82 gnd vdd FILL
XFILL_18_OAI22X1_39 gnd vdd FILL
XFILL_66_DFFSR_93 gnd vdd FILL
XFILL_3_NOR2X1_13 gnd vdd FILL
XFILL_3_NOR2X1_24 gnd vdd FILL
XFILL_44_DFFSR_209 gnd vdd FILL
XFILL_3_NOR2X1_35 gnd vdd FILL
XFILL_3_NOR2X1_46 gnd vdd FILL
XFILL_29_DFFSR_3 gnd vdd FILL
XNAND3X1_70 DFFSR_139/Q BUFX4_92/Y AND2X2_4/A gnd OAI21X1_3/C vdd NAND3X1
XFILL_3_NOR2X1_57 gnd vdd FILL
XFILL_9_DFFSR_40 gnd vdd FILL
XFILL_3_NOR2X1_68 gnd vdd FILL
XFILL_3_NOR2X1_79 gnd vdd FILL
XFILL_86_DFFSR_4 gnd vdd FILL
XFILL_2_CLKBUF1_18 gnd vdd FILL
XNAND3X1_81 DFFSR_25/Q NAND3X1_7/B NOR2X1_38/Y gnd NAND3X1_82/C vdd NAND3X1
XFILL_29_CLKBUF1_2 gnd vdd FILL
XFILL_9_DFFSR_51 gnd vdd FILL
XFILL_2_CLKBUF1_29 gnd vdd FILL
XNAND3X1_92 DFFSR_140/Q BUFX4_92/Y AND2X2_4/A gnd OAI21X1_13/C vdd NAND3X1
XFILL_9_DFFSR_62 gnd vdd FILL
XFILL_71_DFFSR_109 gnd vdd FILL
XFILL_48_DFFSR_208 gnd vdd FILL
XFILL_9_DFFSR_73 gnd vdd FILL
XFILL_7_NOR2X1_12 gnd vdd FILL
XFILL_9_DFFSR_84 gnd vdd FILL
XFILL_7_NOR2X1_23 gnd vdd FILL
XFILL_5_INVX2_1 gnd vdd FILL
XFILL_9_DFFSR_95 gnd vdd FILL
XFILL_48_DFFSR_219 gnd vdd FILL
XFILL_7_NOR2X1_34 gnd vdd FILL
XFILL_35_DFFSR_70 gnd vdd FILL
XFILL_7_NOR2X1_45 gnd vdd FILL
XFILL_35_DFFSR_81 gnd vdd FILL
XFILL_62_4_0 gnd vdd FILL
XFILL_7_NOR2X1_56 gnd vdd FILL
XFILL_35_DFFSR_92 gnd vdd FILL
XFILL_11_OAI22X1_7 gnd vdd FILL
XNOR2X1_70 INVX1_69/Y NOR2X1_86/B gnd NOR3X1_25/C vdd NOR2X1
XFILL_7_NOR2X1_67 gnd vdd FILL
XNOR2X1_81 NOR2X1_81/A NOR2X1_81/B gnd NOR2X1_81/Y vdd NOR2X1
XFILL_7_NOR2X1_78 gnd vdd FILL
XNOR2X1_92 NOR2X1_92/A NOR2X1_92/B gnd NOR2X1_92/Y vdd NOR2X1
XFILL_34_1_2 gnd vdd FILL
XFILL_7_NOR2X1_89 gnd vdd FILL
XFILL_75_DFFSR_108 gnd vdd FILL
XFILL_0_NOR2X1_103 gnd vdd FILL
XFILL_0_NOR2X1_114 gnd vdd FILL
XFILL_75_DFFSR_119 gnd vdd FILL
XFILL_0_NOR2X1_125 gnd vdd FILL
XFILL_11_OAI21X1_19 gnd vdd FILL
XFILL_0_NOR2X1_136 gnd vdd FILL
XFILL_75_DFFSR_80 gnd vdd FILL
XFILL_0_NOR2X1_147 gnd vdd FILL
XFILL_15_OAI22X1_6 gnd vdd FILL
XFILL_75_DFFSR_91 gnd vdd FILL
XFILL_13_DFFSR_9 gnd vdd FILL
XFILL_0_NOR2X1_158 gnd vdd FILL
XFILL_11_2 gnd vdd FILL
XFILL_0_NOR2X1_169 gnd vdd FILL
XFILL_79_DFFSR_107 gnd vdd FILL
XFILL_79_DFFSR_118 gnd vdd FILL
XFILL_10_NAND2X1_40 gnd vdd FILL
XFILL_79_DFFSR_129 gnd vdd FILL
XFILL_10_NAND2X1_51 gnd vdd FILL
XFILL_19_OAI22X1_5 gnd vdd FILL
XFILL_10_NAND2X1_62 gnd vdd FILL
XFILL_10_NAND2X1_73 gnd vdd FILL
XFILL_8_OAI22X1_12 gnd vdd FILL
XFILL_8_OAI22X1_23 gnd vdd FILL
XFILL_10_NAND2X1_84 gnd vdd FILL
XFILL_8_OAI22X1_34 gnd vdd FILL
XFILL_10_NAND2X1_95 gnd vdd FILL
XFILL_8_OAI22X1_45 gnd vdd FILL
XFILL_44_DFFSR_90 gnd vdd FILL
XBUFX2_8 BUFX2_8/A gnd addr[4] vdd BUFX2
XFILL_33_DFFSR_230 gnd vdd FILL
XFILL_33_DFFSR_241 gnd vdd FILL
XFILL_33_DFFSR_252 gnd vdd FILL
XFILL_33_DFFSR_263 gnd vdd FILL
XFILL_33_DFFSR_274 gnd vdd FILL
XFILL_0_MUX2X1_109 gnd vdd FILL
XFILL_5_NOR2X1_203 gnd vdd FILL
XFILL_60_DFFSR_130 gnd vdd FILL
XFILL_37_DFFSR_240 gnd vdd FILL
XFILL_60_DFFSR_141 gnd vdd FILL
XFILL_60_DFFSR_152 gnd vdd FILL
XFILL_37_DFFSR_251 gnd vdd FILL
XFILL_37_DFFSR_262 gnd vdd FILL
XFILL_60_DFFSR_163 gnd vdd FILL
XFILL_60_DFFSR_174 gnd vdd FILL
XNAND2X1_3 OAI21X1_1/A NAND3X1_1/B gnd NAND2X1_3/Y vdd NAND2X1
XFILL_1_OAI21X1_14 gnd vdd FILL
XFILL_37_DFFSR_273 gnd vdd FILL
XFILL_3_MUX2X1_20 gnd vdd FILL
XFILL_60_DFFSR_185 gnd vdd FILL
XFILL_1_OAI21X1_25 gnd vdd FILL
XFILL_3_MUX2X1_31 gnd vdd FILL
XFILL_3_MUX2X1_42 gnd vdd FILL
XFILL_1_OAI21X1_36 gnd vdd FILL
XFILL_19_CLKBUF1_10 gnd vdd FILL
XFILL_60_DFFSR_196 gnd vdd FILL
XFILL_19_CLKBUF1_21 gnd vdd FILL
XFILL_11_DFFSR_209 gnd vdd FILL
XFILL_19_CLKBUF1_32 gnd vdd FILL
XFILL_3_MUX2X1_53 gnd vdd FILL
XFILL_1_OAI21X1_47 gnd vdd FILL
XFILL_64_DFFSR_140 gnd vdd FILL
XFILL_3_MUX2X1_64 gnd vdd FILL
XFILL_3_MUX2X1_75 gnd vdd FILL
XFILL_3_MUX2X1_86 gnd vdd FILL
XFILL_64_DFFSR_151 gnd vdd FILL
XFILL_64_DFFSR_162 gnd vdd FILL
XFILL_3_MUX2X1_97 gnd vdd FILL
XFILL_14_AOI21X1_40 gnd vdd FILL
XFILL_64_DFFSR_173 gnd vdd FILL
XFILL_64_DFFSR_184 gnd vdd FILL
XFILL_14_AOI21X1_51 gnd vdd FILL
XFILL_7_MUX2X1_30 gnd vdd FILL
XFILL_64_DFFSR_195 gnd vdd FILL
XFILL_7_MUX2X1_41 gnd vdd FILL
XFILL_14_AOI21X1_62 gnd vdd FILL
XFILL_53_4_0 gnd vdd FILL
XFILL_15_DFFSR_208 gnd vdd FILL
XFILL_7_MUX2X1_52 gnd vdd FILL
XFILL_14_AOI21X1_73 gnd vdd FILL
XFILL_12_NAND3X1_8 gnd vdd FILL
XFILL_15_DFFSR_219 gnd vdd FILL
XFILL_25_1_2 gnd vdd FILL
XFILL_0_1_2 gnd vdd FILL
XFILL_7_MUX2X1_63 gnd vdd FILL
XFILL_68_DFFSR_150 gnd vdd FILL
XFILL_0_NAND2X1_90 gnd vdd FILL
XFILL_7_MUX2X1_74 gnd vdd FILL
XNOR2X1_160 DFFSR_83/Q NOR2X1_161/B gnd NOR2X1_160/Y vdd NOR2X1
XFILL_7_MUX2X1_85 gnd vdd FILL
XFILL_68_DFFSR_161 gnd vdd FILL
XFILL_7_MUX2X1_96 gnd vdd FILL
XNOR2X1_171 BUFX2_9/A INVX1_136/Y gnd NAND2X1_4/B vdd NOR2X1
XFILL_68_DFFSR_172 gnd vdd FILL
XNOR2X1_182 NOR2X1_7/B NOR2X1_35/B gnd MUX2X1_16/S vdd NOR2X1
XFILL_68_DFFSR_183 gnd vdd FILL
XNOR2X1_193 DFFSR_16/Q NOR2X1_195/B gnd NOR2X1_193/Y vdd NOR2X1
XFILL_68_DFFSR_194 gnd vdd FILL
XFILL_19_DFFSR_207 gnd vdd FILL
XFILL_42_DFFSR_108 gnd vdd FILL
XFILL_42_DFFSR_119 gnd vdd FILL
XFILL_19_DFFSR_218 gnd vdd FILL
XFILL_19_DFFSR_229 gnd vdd FILL
XFILL_46_DFFSR_107 gnd vdd FILL
XAOI21X1_8 BUFX4_87/Y AOI21X1_9/B AOI21X1_8/C gnd DFFSR_103/D vdd AOI21X1
XFILL_46_DFFSR_118 gnd vdd FILL
XFILL_46_DFFSR_129 gnd vdd FILL
XMUX2X1_100 NOR3X1_10/A BUFX4_87/Y NAND2X1_16/Y gnd DFFSR_13/D vdd MUX2X1
XMUX2X1_111 INVX1_153/Y BUFX4_74/Y NAND2X1_23/Y gnd DFFSR_154/D vdd MUX2X1
XMUX2X1_122 BUFX4_83/Y OAI21X1_2/A NOR2X1_136/Y gnd DFFSR_130/D vdd MUX2X1
XMUX2X1_133 INVX1_177/Y BUFX4_77/Y NAND2X1_2/Y gnd DFFSR_123/D vdd MUX2X1
XMUX2X1_144 BUFX4_80/Y OAI21X1_7/A NOR2X1_142/Y gnd DFFSR_107/D vdd MUX2X1
XMUX2X1_155 BUFX4_78/Y INVX1_199/Y NOR2X1_155/Y gnd DFFSR_92/D vdd MUX2X1
XFILL_17_MUX2X1_101 gnd vdd FILL
XFILL_17_MUX2X1_112 gnd vdd FILL
XFILL_17_MUX2X1_123 gnd vdd FILL
XMUX2X1_166 BUFX4_80/Y INVX1_211/Y NOR2X1_164/Y gnd DFFSR_72/D vdd MUX2X1
XFILL_23_MUX2X1_50 gnd vdd FILL
XFILL_23_MUX2X1_61 gnd vdd FILL
XFILL_17_MUX2X1_134 gnd vdd FILL
XMUX2X1_177 BUFX4_74/Y INVX1_222/Y NOR2X1_166/Y gnd DFFSR_65/D vdd MUX2X1
XFILL_17_MUX2X1_145 gnd vdd FILL
XMUX2X1_188 BUFX4_87/Y INVX1_7/Y NOR2X1_169/Y gnd DFFSR_50/D vdd MUX2X1
XFILL_23_MUX2X1_72 gnd vdd FILL
XFILL_23_MUX2X1_83 gnd vdd FILL
XFILL_23_MUX2X1_94 gnd vdd FILL
XFILL_17_MUX2X1_156 gnd vdd FILL
XFILL_9_BUFX2_2 gnd vdd FILL
XFILL_8_2_2 gnd vdd FILL
XFILL_17_MUX2X1_167 gnd vdd FILL
XFILL_17_MUX2X1_178 gnd vdd FILL
XFILL_17_MUX2X1_189 gnd vdd FILL
XINVX1_40 INVX1_40/A gnd INVX1_40/Y vdd INVX1
XINVX1_51 INVX1_51/A gnd INVX1_51/Y vdd INVX1
XFILL_30_DFFSR_3 gnd vdd FILL
XINVX1_62 INVX1_62/A gnd INVX1_62/Y vdd INVX1
XINVX1_73 INVX1_73/A gnd INVX1_73/Y vdd INVX1
XINVX1_84 INVX1_84/A gnd INVX1_84/Y vdd INVX1
XINVX1_95 INVX1_95/A gnd INVX1_95/Y vdd INVX1
XFILL_68_DFFSR_1 gnd vdd FILL
XFILL_3_INVX1_17 gnd vdd FILL
XFILL_3_INVX1_28 gnd vdd FILL
XFILL_31_DFFSR_140 gnd vdd FILL
XFILL_31_DFFSR_151 gnd vdd FILL
XFILL_3_INVX1_39 gnd vdd FILL
XFILL_31_DFFSR_162 gnd vdd FILL
XFILL_44_4_0 gnd vdd FILL
XFILL_31_DFFSR_173 gnd vdd FILL
XFILL_16_1_2 gnd vdd FILL
XFILL_31_DFFSR_184 gnd vdd FILL
XFILL_31_DFFSR_195 gnd vdd FILL
XFILL_35_DFFSR_150 gnd vdd FILL
XFILL_35_DFFSR_161 gnd vdd FILL
XFILL_35_DFFSR_172 gnd vdd FILL
XFILL_35_DFFSR_183 gnd vdd FILL
XFILL_35_DFFSR_194 gnd vdd FILL
XFILL_1_BUFX4_15 gnd vdd FILL
XFILL_1_BUFX4_26 gnd vdd FILL
XFILL_52_DFFSR_7 gnd vdd FILL
XFILL_7_MUX2X1_140 gnd vdd FILL
XFILL_1_BUFX4_37 gnd vdd FILL
XFILL_1_BUFX4_48 gnd vdd FILL
XFILL_7_MUX2X1_151 gnd vdd FILL
XFILL_18_DFFSR_19 gnd vdd FILL
XFILL_7_MUX2X1_162 gnd vdd FILL
XFILL_1_BUFX4_59 gnd vdd FILL
XFILL_39_DFFSR_160 gnd vdd FILL
XFILL_7_MUX2X1_173 gnd vdd FILL
XFILL_39_DFFSR_171 gnd vdd FILL
XFILL_7_MUX2X1_184 gnd vdd FILL
XFILL_39_DFFSR_182 gnd vdd FILL
XFILL_39_DFFSR_193 gnd vdd FILL
XFILL_13_DFFSR_107 gnd vdd FILL
XFILL_13_DFFSR_118 gnd vdd FILL
XFILL_31_NOR3X1_40 gnd vdd FILL
XFILL_31_NOR3X1_51 gnd vdd FILL
XFILL_13_DFFSR_129 gnd vdd FILL
XFILL_58_DFFSR_18 gnd vdd FILL
XNOR2X1_6 NOR2X1_6/A NOR2X1_6/B gnd NOR2X1_6/Y vdd NOR2X1
XFILL_58_DFFSR_29 gnd vdd FILL
XFILL_81_DFFSR_240 gnd vdd FILL
XFILL_81_DFFSR_251 gnd vdd FILL
XFILL_81_DFFSR_262 gnd vdd FILL
XFILL_17_DFFSR_106 gnd vdd FILL
XFILL_81_DFFSR_273 gnd vdd FILL
XFILL_17_DFFSR_117 gnd vdd FILL
XFILL_17_DFFSR_128 gnd vdd FILL
XFILL_17_DFFSR_139 gnd vdd FILL
XFILL_12_AOI21X1_2 gnd vdd FILL
XFILL_85_DFFSR_250 gnd vdd FILL
XFILL_85_DFFSR_261 gnd vdd FILL
XFILL_27_DFFSR_17 gnd vdd FILL
XFILL_85_DFFSR_272 gnd vdd FILL
XFILL_27_DFFSR_28 gnd vdd FILL
XFILL_66_3 gnd vdd FILL
XFILL_27_DFFSR_39 gnd vdd FILL
XFILL_66_0_2 gnd vdd FILL
XFILL_59_2 gnd vdd FILL
XFILL_13_NOR3X1_18 gnd vdd FILL
XFILL_67_DFFSR_16 gnd vdd FILL
XFILL_67_DFFSR_27 gnd vdd FILL
XFILL_8_NAND3X1_130 gnd vdd FILL
XFILL_13_NOR3X1_29 gnd vdd FILL
XFILL_67_DFFSR_38 gnd vdd FILL
XFILL_35_4_0 gnd vdd FILL
XFILL_63_DFFSR_207 gnd vdd FILL
XFILL_67_DFFSR_49 gnd vdd FILL
XFILL_63_DFFSR_218 gnd vdd FILL
XFILL_63_DFFSR_229 gnd vdd FILL
XFILL_17_NOR3X1_17 gnd vdd FILL
XFILL_17_NOR3X1_28 gnd vdd FILL
XFILL_17_NOR3X1_39 gnd vdd FILL
XFILL_67_DFFSR_206 gnd vdd FILL
XFILL_67_DFFSR_217 gnd vdd FILL
XFILL_36_DFFSR_15 gnd vdd FILL
XFILL_36_DFFSR_26 gnd vdd FILL
XFILL_67_DFFSR_228 gnd vdd FILL
XFILL_36_DFFSR_37 gnd vdd FILL
XFILL_67_DFFSR_239 gnd vdd FILL
XFILL_36_DFFSR_48 gnd vdd FILL
XFILL_36_DFFSR_59 gnd vdd FILL
XAOI21X1_16 MUX2X1_2/A NOR2X1_153/B NOR2X1_153/Y gnd DFFSR_102/D vdd AOI21X1
XAOI21X1_27 MUX2X1_66/A NOR2X1_181/B NOR2X1_181/Y gnd DFFSR_31/D vdd AOI21X1
XFILL_76_DFFSR_14 gnd vdd FILL
XAOI21X1_38 BUFX4_99/Y NOR2X1_195/B NOR2X1_195/Y gnd DFFSR_18/D vdd AOI21X1
XAOI21X1_49 BUFX4_97/Y NOR2X1_6/B NOR2X1_6/Y gnd DFFSR_274/D vdd AOI21X1
XFILL_76_DFFSR_25 gnd vdd FILL
XFILL_76_DFFSR_36 gnd vdd FILL
XFILL_3_NAND2X1_12 gnd vdd FILL
XFILL_76_DFFSR_47 gnd vdd FILL
XFILL_76_DFFSR_58 gnd vdd FILL
XFILL_19_MUX2X1_4 gnd vdd FILL
XFILL_3_NAND2X1_23 gnd vdd FILL
XFILL_76_DFFSR_69 gnd vdd FILL
XFILL_3_NAND2X1_34 gnd vdd FILL
XFILL_3_NAND2X1_45 gnd vdd FILL
XFILL_3_NAND2X1_56 gnd vdd FILL
XFILL_3_NAND2X1_67 gnd vdd FILL
XFILL_3_NAND2X1_78 gnd vdd FILL
XFILL_0_AND2X2_2 gnd vdd FILL
XFILL_3_NAND2X1_89 gnd vdd FILL
XFILL_45_DFFSR_13 gnd vdd FILL
XFILL_45_DFFSR_24 gnd vdd FILL
XFILL_45_DFFSR_35 gnd vdd FILL
XFILL_45_DFFSR_46 gnd vdd FILL
XFILL_45_DFFSR_57 gnd vdd FILL
XFILL_45_DFFSR_68 gnd vdd FILL
XFILL_45_DFFSR_79 gnd vdd FILL
XFILL_85_DFFSR_12 gnd vdd FILL
XFILL_52_DFFSR_250 gnd vdd FILL
XFILL_85_DFFSR_23 gnd vdd FILL
XFILL_52_DFFSR_261 gnd vdd FILL
XFILL_57_0_2 gnd vdd FILL
XFILL_52_DFFSR_272 gnd vdd FILL
XFILL_85_DFFSR_34 gnd vdd FILL
XFILL_85_DFFSR_45 gnd vdd FILL
XFILL_29_CLKBUF1_11 gnd vdd FILL
XFILL_85_DFFSR_56 gnd vdd FILL
XFILL_14_DFFSR_12 gnd vdd FILL
XFILL_29_CLKBUF1_22 gnd vdd FILL
XFILL_85_DFFSR_67 gnd vdd FILL
XFILL_14_DFFSR_23 gnd vdd FILL
XFILL_85_DFFSR_78 gnd vdd FILL
XFILL_29_CLKBUF1_33 gnd vdd FILL
XFILL_14_DFFSR_34 gnd vdd FILL
XFILL_85_DFFSR_89 gnd vdd FILL
XFILL_14_DFFSR_45 gnd vdd FILL
XFILL_14_DFFSR_56 gnd vdd FILL
XFILL_3_AOI22X1_10 gnd vdd FILL
XFILL_14_DFFSR_67 gnd vdd FILL
XFILL_1_4_0 gnd vdd FILL
XFILL_56_DFFSR_260 gnd vdd FILL
XFILL_26_4_0 gnd vdd FILL
XFILL_14_DFFSR_78 gnd vdd FILL
XFILL_11_CLKBUF1_1 gnd vdd FILL
XFILL_56_DFFSR_271 gnd vdd FILL
XFILL_14_DFFSR_89 gnd vdd FILL
XFILL_54_DFFSR_11 gnd vdd FILL
XFILL_30_DFFSR_207 gnd vdd FILL
XFILL_7_AOI21X1_12 gnd vdd FILL
XFILL_54_DFFSR_22 gnd vdd FILL
XFILL_30_DFFSR_218 gnd vdd FILL
XFILL_54_DFFSR_33 gnd vdd FILL
XOAI22X1_13 INVX1_198/Y OAI22X1_49/B INVX1_202/Y OAI22X1_49/D gnd NOR2X1_64/A vdd
+ OAI22X1
XFILL_25_NOR3X1_8 gnd vdd FILL
XFILL_30_DFFSR_229 gnd vdd FILL
XOAI22X1_24 INVX1_199/Y OAI22X1_49/B INVX1_203/Y OAI22X1_49/D gnd NOR2X1_83/A vdd
+ OAI22X1
XFILL_7_AOI21X1_23 gnd vdd FILL
XFILL_7_AOI21X1_34 gnd vdd FILL
XOAI22X1_35 INVX1_75/Y OAI22X1_1/B INVX1_80/Y OAI22X1_1/D gnd NOR3X1_38/C vdd OAI22X1
XFILL_54_DFFSR_44 gnd vdd FILL
XFILL_7_AOI21X1_45 gnd vdd FILL
XFILL_54_DFFSR_55 gnd vdd FILL
XOAI22X1_46 INVX1_6/Y OAI22X1_5/B INVX1_11/Y OAI22X1_5/D gnd OAI22X1_46/Y vdd OAI22X1
XFILL_83_DFFSR_160 gnd vdd FILL
XFILL_54_DFFSR_66 gnd vdd FILL
XFILL_7_AOI21X1_56 gnd vdd FILL
XFILL_54_DFFSR_77 gnd vdd FILL
XFILL_17_OAI22X1_14 gnd vdd FILL
XFILL_83_DFFSR_171 gnd vdd FILL
XFILL_7_AOI21X1_67 gnd vdd FILL
XFILL_54_DFFSR_88 gnd vdd FILL
XFILL_17_OAI22X1_25 gnd vdd FILL
XFILL_83_DFFSR_182 gnd vdd FILL
XFILL_7_AOI21X1_78 gnd vdd FILL
XFILL_83_DFFSR_193 gnd vdd FILL
XFILL_17_OAI22X1_36 gnd vdd FILL
XFILL_34_DFFSR_206 gnd vdd FILL
XFILL_54_DFFSR_99 gnd vdd FILL
XFILL_17_OAI22X1_47 gnd vdd FILL
XFILL_34_DFFSR_217 gnd vdd FILL
XFILL_3_DFFSR_230 gnd vdd FILL
XFILL_3_DFFSR_241 gnd vdd FILL
XFILL_34_DFFSR_228 gnd vdd FILL
XFILL_34_DFFSR_4 gnd vdd FILL
XFILL_34_DFFSR_239 gnd vdd FILL
XFILL_3_DFFSR_252 gnd vdd FILL
XFILL_23_DFFSR_10 gnd vdd FILL
XFILL_3_DFFSR_263 gnd vdd FILL
XFILL_23_DFFSR_21 gnd vdd FILL
XFILL_1_CLKBUF1_15 gnd vdd FILL
XFILL_3_DFFSR_274 gnd vdd FILL
XFILL_87_DFFSR_170 gnd vdd FILL
XFILL_23_DFFSR_32 gnd vdd FILL
XFILL_23_DFFSR_43 gnd vdd FILL
XFILL_0_MUX2X1_19 gnd vdd FILL
XFILL_1_CLKBUF1_26 gnd vdd FILL
XFILL_87_DFFSR_181 gnd vdd FILL
XFILL_87_DFFSR_192 gnd vdd FILL
XFILL_1_CLKBUF1_37 gnd vdd FILL
XFILL_61_DFFSR_106 gnd vdd FILL
XFILL_38_DFFSR_205 gnd vdd FILL
XFILL_23_DFFSR_54 gnd vdd FILL
XFILL_38_DFFSR_216 gnd vdd FILL
XFILL_23_DFFSR_65 gnd vdd FILL
XFILL_61_DFFSR_117 gnd vdd FILL
XFILL_23_DFFSR_76 gnd vdd FILL
XFILL_61_DFFSR_128 gnd vdd FILL
XFILL_38_DFFSR_227 gnd vdd FILL
XFILL_23_DFFSR_87 gnd vdd FILL
XFILL_7_DFFSR_240 gnd vdd FILL
XFILL_23_DFFSR_98 gnd vdd FILL
XFILL_7_DFFSR_251 gnd vdd FILL
XFILL_38_DFFSR_238 gnd vdd FILL
XFILL_61_DFFSR_139 gnd vdd FILL
XFILL_8_NOR3X1_9 gnd vdd FILL
XFILL_38_DFFSR_249 gnd vdd FILL
XFILL_7_DFFSR_262 gnd vdd FILL
XFILL_63_DFFSR_20 gnd vdd FILL
XFILL_7_DFFSR_273 gnd vdd FILL
XFILL_63_DFFSR_31 gnd vdd FILL
XFILL_4_MUX2X1_18 gnd vdd FILL
XFILL_63_DFFSR_42 gnd vdd FILL
XFILL_4_MUX2X1_29 gnd vdd FILL
XFILL_63_DFFSR_53 gnd vdd FILL
XFILL_65_DFFSR_105 gnd vdd FILL
XFILL_10_OAI21X1_16 gnd vdd FILL
XFILL_65_DFFSR_116 gnd vdd FILL
XFILL_63_DFFSR_64 gnd vdd FILL
XFILL_65_DFFSR_127 gnd vdd FILL
XFILL_9_5_0 gnd vdd FILL
XFILL_63_DFFSR_75 gnd vdd FILL
XFILL_65_DFFSR_138 gnd vdd FILL
XFILL_10_OAI21X1_27 gnd vdd FILL
XFILL_63_DFFSR_86 gnd vdd FILL
XFILL_10_OAI21X1_38 gnd vdd FILL
XFILL_63_DFFSR_97 gnd vdd FILL
XFILL_65_DFFSR_149 gnd vdd FILL
XFILL_10_OAI21X1_49 gnd vdd FILL
XFILL_6_DFFSR_11 gnd vdd FILL
XFILL_6_DFFSR_22 gnd vdd FILL
XFILL_8_MUX2X1_17 gnd vdd FILL
XFILL_6_DFFSR_33 gnd vdd FILL
XFILL_8_MUX2X1_28 gnd vdd FILL
XFILL_69_DFFSR_104 gnd vdd FILL
XFILL_8_MUX2X1_39 gnd vdd FILL
XFILL_6_DFFSR_44 gnd vdd FILL
XFILL_56_DFFSR_8 gnd vdd FILL
XFILL_69_DFFSR_115 gnd vdd FILL
XFILL_6_DFFSR_55 gnd vdd FILL
XFILL_69_DFFSR_126 gnd vdd FILL
XFILL_32_DFFSR_30 gnd vdd FILL
XFILL_69_DFFSR_137 gnd vdd FILL
XFILL_48_0_2 gnd vdd FILL
XFILL_6_DFFSR_66 gnd vdd FILL
XFILL_0_AOI22X1_2 gnd vdd FILL
XFILL_32_DFFSR_41 gnd vdd FILL
XFILL_6_DFFSR_77 gnd vdd FILL
XFILL_69_DFFSR_148 gnd vdd FILL
XFILL_32_DFFSR_52 gnd vdd FILL
XFILL_32_DFFSR_63 gnd vdd FILL
XFILL_12_OAI21X1_5 gnd vdd FILL
XFILL_6_DFFSR_88 gnd vdd FILL
XFILL_6_DFFSR_99 gnd vdd FILL
XFILL_7_OAI22X1_20 gnd vdd FILL
XFILL_69_DFFSR_159 gnd vdd FILL
XFILL_7_OAI22X1_31 gnd vdd FILL
XFILL_32_DFFSR_74 gnd vdd FILL
XFILL_7_OAI22X1_42 gnd vdd FILL
XFILL_32_DFFSR_85 gnd vdd FILL
XFILL_32_DFFSR_96 gnd vdd FILL
XFILL_0_INVX1_201 gnd vdd FILL
XFILL_0_INVX1_212 gnd vdd FILL
XFILL_0_INVX1_223 gnd vdd FILL
XFILL_17_4_0 gnd vdd FILL
XFILL_72_DFFSR_40 gnd vdd FILL
XFILL_4_AOI22X1_1 gnd vdd FILL
XFILL_72_DFFSR_51 gnd vdd FILL
XFILL_72_DFFSR_62 gnd vdd FILL
XFILL_72_DFFSR_73 gnd vdd FILL
XFILL_23_DFFSR_260 gnd vdd FILL
XFILL_72_DFFSR_84 gnd vdd FILL
XFILL_60_7_1 gnd vdd FILL
XFILL_72_DFFSR_95 gnd vdd FILL
XFILL_23_DFFSR_271 gnd vdd FILL
XFILL_4_INVX1_200 gnd vdd FILL
XFILL_20_MUX2X1_16 gnd vdd FILL
XFILL_4_INVX1_211 gnd vdd FILL
XFILL_20_MUX2X1_27 gnd vdd FILL
XFILL_4_NOR2X1_200 gnd vdd FILL
XFILL_20_MUX2X1_38 gnd vdd FILL
XFILL_4_INVX1_222 gnd vdd FILL
XFILL_20_MUX2X1_49 gnd vdd FILL
XFILL_50_DFFSR_160 gnd vdd FILL
XFILL_12_NOR3X1_3 gnd vdd FILL
XFILL_27_DFFSR_270 gnd vdd FILL
XFILL_50_DFFSR_171 gnd vdd FILL
XFILL_0_OAI21X1_11 gnd vdd FILL
XFILL_50_DFFSR_182 gnd vdd FILL
XFILL_41_DFFSR_50 gnd vdd FILL
XFILL_50_DFFSR_193 gnd vdd FILL
XFILL_0_OAI21X1_22 gnd vdd FILL
XFILL_41_DFFSR_61 gnd vdd FILL
XFILL_0_OAI21X1_33 gnd vdd FILL
XFILL_41_DFFSR_72 gnd vdd FILL
XFILL_41_DFFSR_83 gnd vdd FILL
XFILL_0_OAI21X1_44 gnd vdd FILL
XFILL_41_DFFSR_94 gnd vdd FILL
XFILL_18_CLKBUF1_40 gnd vdd FILL
XFILL_54_DFFSR_170 gnd vdd FILL
XFILL_54_DFFSR_181 gnd vdd FILL
XFILL_81_DFFSR_60 gnd vdd FILL
XFILL_54_DFFSR_192 gnd vdd FILL
XFILL_81_DFFSR_71 gnd vdd FILL
XFILL_81_DFFSR_82 gnd vdd FILL
XFILL_13_AOI21X1_70 gnd vdd FILL
XFILL_13_AOI21X1_81 gnd vdd FILL
XFILL_81_DFFSR_93 gnd vdd FILL
XFILL_10_DFFSR_60 gnd vdd FILL
XFILL_10_DFFSR_71 gnd vdd FILL
XFILL_10_DFFSR_82 gnd vdd FILL
XFILL_10_DFFSR_93 gnd vdd FILL
XFILL_58_DFFSR_180 gnd vdd FILL
XFILL_58_DFFSR_191 gnd vdd FILL
XFILL_32_DFFSR_105 gnd vdd FILL
XFILL_32_DFFSR_116 gnd vdd FILL
XFILL_21_NOR3X1_1 gnd vdd FILL
XFILL_1_DFFSR_140 gnd vdd FILL
XFILL_32_DFFSR_127 gnd vdd FILL
XFILL_32_DFFSR_138 gnd vdd FILL
XFILL_1_DFFSR_151 gnd vdd FILL
XFILL_1_DFFSR_162 gnd vdd FILL
XFILL_32_DFFSR_149 gnd vdd FILL
XFILL_50_DFFSR_70 gnd vdd FILL
XFILL_21_12 gnd vdd FILL
XFILL_1_DFFSR_173 gnd vdd FILL
XFILL_50_DFFSR_81 gnd vdd FILL
XFILL_1_DFFSR_184 gnd vdd FILL
XFILL_50_DFFSR_92 gnd vdd FILL
XFILL_39_0_2 gnd vdd FILL
XFILL_1_DFFSR_195 gnd vdd FILL
XFILL_36_DFFSR_104 gnd vdd FILL
XFILL_36_DFFSR_115 gnd vdd FILL
XFILL_36_DFFSR_126 gnd vdd FILL
XFILL_36_DFFSR_137 gnd vdd FILL
XFILL_5_DFFSR_150 gnd vdd FILL
XFILL_36_DFFSR_148 gnd vdd FILL
XFILL_5_DFFSR_161 gnd vdd FILL
XFILL_5_DFFSR_172 gnd vdd FILL
XFILL_36_DFFSR_159 gnd vdd FILL
XFILL_5_DFFSR_183 gnd vdd FILL
XFILL_5_DFFSR_194 gnd vdd FILL
XFILL_9_NAND3X1_120 gnd vdd FILL
XFILL_9_NAND3X1_131 gnd vdd FILL
XFILL_4_NOR3X1_2 gnd vdd FILL
XFILL_9_DFFSR_160 gnd vdd FILL
XFILL_16_MUX2X1_120 gnd vdd FILL
XFILL_51_7_1 gnd vdd FILL
XFILL_16_MUX2X1_131 gnd vdd FILL
XFILL_16_MUX2X1_142 gnd vdd FILL
XFILL_9_DFFSR_171 gnd vdd FILL
XFILL_13_MUX2X1_80 gnd vdd FILL
XFILL_16_MUX2X1_153 gnd vdd FILL
XFILL_9_DFFSR_182 gnd vdd FILL
XFILL_13_MUX2X1_91 gnd vdd FILL
XFILL_50_2_0 gnd vdd FILL
XFILL_9_DFFSR_193 gnd vdd FILL
XFILL_16_MUX2X1_164 gnd vdd FILL
XFILL_16_MUX2X1_175 gnd vdd FILL
XFILL_1_NOR3X1_40 gnd vdd FILL
XFILL_1_NOR3X1_51 gnd vdd FILL
XFILL_16_MUX2X1_186 gnd vdd FILL
XFILL_82_DFFSR_205 gnd vdd FILL
XFILL_82_DFFSR_216 gnd vdd FILL
XFILL_82_DFFSR_227 gnd vdd FILL
XFILL_3_DFFSR_3 gnd vdd FILL
XFILL_82_DFFSR_238 gnd vdd FILL
XFILL_82_DFFSR_249 gnd vdd FILL
XFILL_17_MUX2X1_90 gnd vdd FILL
XFILL_16_DFFSR_1 gnd vdd FILL
XFILL_5_NOR3X1_50 gnd vdd FILL
XFILL_73_DFFSR_2 gnd vdd FILL
XFILL_2_DFFSR_70 gnd vdd FILL
XFILL_86_DFFSR_204 gnd vdd FILL
XFILL_86_DFFSR_215 gnd vdd FILL
XFILL_2_DFFSR_81 gnd vdd FILL
XFILL_2_DFFSR_92 gnd vdd FILL
XFILL_86_DFFSR_226 gnd vdd FILL
XFILL_86_DFFSR_237 gnd vdd FILL
XFILL_86_DFFSR_248 gnd vdd FILL
XFILL_21_DFFSR_170 gnd vdd FILL
XFILL_86_DFFSR_259 gnd vdd FILL
XFILL_21_DFFSR_181 gnd vdd FILL
XFILL_2_INVX1_110 gnd vdd FILL
XFILL_21_DFFSR_192 gnd vdd FILL
XFILL_11_BUFX2_7 gnd vdd FILL
XFILL_2_INVX1_121 gnd vdd FILL
XFILL_2_INVX1_132 gnd vdd FILL
XFILL_2_INVX1_143 gnd vdd FILL
XFILL_2_INVX1_154 gnd vdd FILL
XFILL_2_INVX1_165 gnd vdd FILL
XFILL_2_INVX1_176 gnd vdd FILL
XFILL_2_INVX1_187 gnd vdd FILL
XFILL_25_DFFSR_180 gnd vdd FILL
XFILL_2_INVX1_198 gnd vdd FILL
XFILL_25_DFFSR_191 gnd vdd FILL
XFILL_6_INVX1_120 gnd vdd FILL
XFILL_6_INVX1_131 gnd vdd FILL
XFILL_58_3_0 gnd vdd FILL
XFILL_6_INVX1_142 gnd vdd FILL
XFILL_6_INVX1_153 gnd vdd FILL
XFILL_38_DFFSR_5 gnd vdd FILL
XFILL_5_0_2 gnd vdd FILL
XFILL_6_INVX1_164 gnd vdd FILL
XFILL_6_MUX2X1_170 gnd vdd FILL
XFILL_6_INVX1_175 gnd vdd FILL
XFILL_6_INVX1_186 gnd vdd FILL
XFILL_6_INVX1_197 gnd vdd FILL
XFILL_6_MUX2X1_181 gnd vdd FILL
XFILL_29_DFFSR_190 gnd vdd FILL
XFILL_6_MUX2X1_192 gnd vdd FILL
XFILL_0_OAI22X1_5 gnd vdd FILL
XFILL_71_DFFSR_270 gnd vdd FILL
XFILL_42_7_1 gnd vdd FILL
XFILL_41_2_0 gnd vdd FILL
XFILL_4_OAI22X1_4 gnd vdd FILL
XFILL_10_BUFX4_1 gnd vdd FILL
XFILL_8_OAI22X1_3 gnd vdd FILL
XFILL_53_DFFSR_204 gnd vdd FILL
XFILL_53_DFFSR_215 gnd vdd FILL
XFILL_53_DFFSR_226 gnd vdd FILL
XFILL_53_DFFSR_237 gnd vdd FILL
XFILL_9_NAND3X1_40 gnd vdd FILL
XFILL_53_DFFSR_248 gnd vdd FILL
XFILL_9_NAND3X1_51 gnd vdd FILL
XFILL_53_DFFSR_259 gnd vdd FILL
XFILL_9_NAND3X1_62 gnd vdd FILL
XFILL_15_BUFX4_20 gnd vdd FILL
XFILL_9_NAND3X1_73 gnd vdd FILL
XFILL_9_NAND3X1_84 gnd vdd FILL
XFILL_80_DFFSR_104 gnd vdd FILL
XFILL_15_BUFX4_31 gnd vdd FILL
XFILL_9_NAND3X1_95 gnd vdd FILL
XFILL_57_DFFSR_203 gnd vdd FILL
XFILL_15_BUFX4_42 gnd vdd FILL
XFILL_80_DFFSR_115 gnd vdd FILL
XFILL_57_DFFSR_214 gnd vdd FILL
XFILL_15_BUFX4_53 gnd vdd FILL
XFILL_80_DFFSR_126 gnd vdd FILL
XFILL_1_5 gnd vdd FILL
XFILL_15_BUFX4_64 gnd vdd FILL
XFILL_80_DFFSR_137 gnd vdd FILL
XFILL_57_DFFSR_225 gnd vdd FILL
XFILL_57_DFFSR_236 gnd vdd FILL
XFILL_80_DFFSR_148 gnd vdd FILL
XFILL_57_DFFSR_247 gnd vdd FILL
XFILL_15_BUFX4_75 gnd vdd FILL
XFILL_57_DFFSR_258 gnd vdd FILL
XFILL_80_DFFSR_159 gnd vdd FILL
XFILL_15_BUFX4_86 gnd vdd FILL
XFILL_15_BUFX4_97 gnd vdd FILL
XFILL_57_DFFSR_269 gnd vdd FILL
XFILL_49_3_0 gnd vdd FILL
XFILL_0_DFFSR_207 gnd vdd FILL
XFILL_84_DFFSR_103 gnd vdd FILL
XFILL_84_DFFSR_114 gnd vdd FILL
XFILL_0_DFFSR_218 gnd vdd FILL
XFILL_0_DFFSR_229 gnd vdd FILL
XFILL_84_DFFSR_125 gnd vdd FILL
XFILL_84_DFFSR_136 gnd vdd FILL
XFILL_84_DFFSR_147 gnd vdd FILL
XFILL_84_DFFSR_158 gnd vdd FILL
XFILL_43_5 gnd vdd FILL
XFILL_84_DFFSR_169 gnd vdd FILL
XFILL_2_NAND2X1_20 gnd vdd FILL
XFILL_16_CLKBUF1_9 gnd vdd FILL
XFILL_10_INVX4_1 gnd vdd FILL
XFILL_2_NAND2X1_31 gnd vdd FILL
XFILL_4_DFFSR_206 gnd vdd FILL
XFILL_2_NAND2X1_42 gnd vdd FILL
XFILL_2_NAND2X1_53 gnd vdd FILL
XFILL_1_NAND3X1_6 gnd vdd FILL
XFILL_4_DFFSR_217 gnd vdd FILL
XFILL_2_NAND2X1_64 gnd vdd FILL
XFILL_4_DFFSR_228 gnd vdd FILL
XFILL_0_INVX8_1 gnd vdd FILL
XFILL_4_DFFSR_239 gnd vdd FILL
XFILL_2_NAND2X1_75 gnd vdd FILL
XFILL_2_NAND2X1_86 gnd vdd FILL
XFILL_33_7_1 gnd vdd FILL
XFILL_33_DFFSR_19 gnd vdd FILL
XFILL_12_BUFX4_104 gnd vdd FILL
XFILL_32_2_0 gnd vdd FILL
XFILL_8_DFFSR_205 gnd vdd FILL
XFILL_8_DFFSR_216 gnd vdd FILL
XFILL_5_NAND3X1_5 gnd vdd FILL
XFILL_10_CLKBUF1_17 gnd vdd FILL
XFILL_10_CLKBUF1_28 gnd vdd FILL
XFILL_8_DFFSR_227 gnd vdd FILL
XFILL_10_CLKBUF1_39 gnd vdd FILL
XFILL_8_DFFSR_238 gnd vdd FILL
XFILL_8_DFFSR_249 gnd vdd FILL
XFILL_73_DFFSR_18 gnd vdd FILL
XFILL_73_DFFSR_29 gnd vdd FILL
XFILL_16_MUX2X1_8 gnd vdd FILL
XFILL_9_NAND3X1_4 gnd vdd FILL
XFILL_16_12 gnd vdd FILL
XFILL_28_CLKBUF1_30 gnd vdd FILL
XFILL_28_CLKBUF1_41 gnd vdd FILL
XFILL_7_BUFX4_30 gnd vdd FILL
XFILL_7_BUFX4_41 gnd vdd FILL
XFILL_7_BUFX4_52 gnd vdd FILL
XFILL_7_BUFX4_63 gnd vdd FILL
XFILL_42_DFFSR_17 gnd vdd FILL
XFILL_7_BUFX4_74 gnd vdd FILL
XFILL_20_DFFSR_204 gnd vdd FILL
XFILL_7_BUFX4_85 gnd vdd FILL
XFILL_42_DFFSR_28 gnd vdd FILL
XFILL_20_DFFSR_215 gnd vdd FILL
XFILL_6_AOI21X1_20 gnd vdd FILL
XFILL_42_DFFSR_39 gnd vdd FILL
XFILL_19_MUX2X1_108 gnd vdd FILL
XFILL_10_NOR2X1_17 gnd vdd FILL
XFILL_19_MUX2X1_119 gnd vdd FILL
XFILL_7_BUFX4_96 gnd vdd FILL
XFILL_20_DFFSR_226 gnd vdd FILL
XFILL_10_NOR2X1_28 gnd vdd FILL
XFILL_20_DFFSR_237 gnd vdd FILL
XFILL_6_AOI21X1_31 gnd vdd FILL
XFILL_10_NOR2X1_39 gnd vdd FILL
XFILL_6_AOI21X1_42 gnd vdd FILL
XFILL_20_DFFSR_248 gnd vdd FILL
XFILL_6_AOI21X1_53 gnd vdd FILL
XFILL_20_DFFSR_259 gnd vdd FILL
XFILL_16_OAI22X1_11 gnd vdd FILL
XFILL_6_AOI21X1_64 gnd vdd FILL
XFILL_16_OAI22X1_22 gnd vdd FILL
XFILL_73_DFFSR_190 gnd vdd FILL
XFILL_82_DFFSR_16 gnd vdd FILL
XFILL_6_AOI21X1_75 gnd vdd FILL
XFILL_16_OAI22X1_33 gnd vdd FILL
XFILL_16_OAI22X1_44 gnd vdd FILL
XFILL_24_DFFSR_203 gnd vdd FILL
XFILL_82_DFFSR_27 gnd vdd FILL
XFILL_24_DFFSR_214 gnd vdd FILL
XFILL_82_DFFSR_38 gnd vdd FILL
XFILL_82_DFFSR_49 gnd vdd FILL
XFILL_24_DFFSR_225 gnd vdd FILL
XFILL_7_DFFSR_4 gnd vdd FILL
XFILL_11_DFFSR_16 gnd vdd FILL
XFILL_24_DFFSR_236 gnd vdd FILL
XFILL_9_NOR2X1_130 gnd vdd FILL
XFILL_9_NOR2X1_141 gnd vdd FILL
XFILL_24_DFFSR_247 gnd vdd FILL
XFILL_11_DFFSR_27 gnd vdd FILL
XFILL_0_CLKBUF1_12 gnd vdd FILL
XFILL_24_DFFSR_258 gnd vdd FILL
XFILL_9_NOR2X1_152 gnd vdd FILL
XFILL_0_CLKBUF1_23 gnd vdd FILL
XFILL_11_DFFSR_38 gnd vdd FILL
XFILL_24_DFFSR_269 gnd vdd FILL
XFILL_11_DFFSR_49 gnd vdd FILL
XFILL_9_NOR2X1_163 gnd vdd FILL
XFILL_77_DFFSR_3 gnd vdd FILL
XFILL_0_CLKBUF1_34 gnd vdd FILL
XFILL_5_INVX1_209 gnd vdd FILL
XFILL_9_NOR2X1_174 gnd vdd FILL
XFILL_28_DFFSR_202 gnd vdd FILL
XFILL_51_DFFSR_103 gnd vdd FILL
XFILL_9_NOR2X1_185 gnd vdd FILL
XFILL_9_NOR2X1_9 gnd vdd FILL
XFILL_28_DFFSR_213 gnd vdd FILL
XFILL_51_DFFSR_114 gnd vdd FILL
XFILL_9_NOR2X1_196 gnd vdd FILL
XFILL_51_DFFSR_125 gnd vdd FILL
XFILL_51_DFFSR_136 gnd vdd FILL
XFILL_9_AOI22X1_9 gnd vdd FILL
XFILL_28_DFFSR_224 gnd vdd FILL
XFILL_28_DFFSR_235 gnd vdd FILL
XFILL_51_DFFSR_15 gnd vdd FILL
XFILL_51_DFFSR_26 gnd vdd FILL
XFILL_28_DFFSR_246 gnd vdd FILL
XFILL_51_DFFSR_147 gnd vdd FILL
XFILL_51_DFFSR_158 gnd vdd FILL
XFILL_51_DFFSR_37 gnd vdd FILL
XFILL_28_DFFSR_257 gnd vdd FILL
XFILL_28_DFFSR_268 gnd vdd FILL
XFILL_51_DFFSR_169 gnd vdd FILL
XFILL_51_DFFSR_48 gnd vdd FILL
XFILL_51_DFFSR_59 gnd vdd FILL
XFILL_55_DFFSR_102 gnd vdd FILL
XFILL_24_7_1 gnd vdd FILL
XFILL_55_DFFSR_113 gnd vdd FILL
XFILL_55_DFFSR_124 gnd vdd FILL
XFILL_23_2_0 gnd vdd FILL
XFILL_55_DFFSR_135 gnd vdd FILL
XFILL_55_DFFSR_146 gnd vdd FILL
XFILL_8_MUX2X1_7 gnd vdd FILL
XFILL_55_DFFSR_157 gnd vdd FILL
XFILL_55_DFFSR_168 gnd vdd FILL
XFILL_55_DFFSR_179 gnd vdd FILL
XFILL_9_MUX2X1_103 gnd vdd FILL
XFILL_59_DFFSR_101 gnd vdd FILL
XFILL_20_DFFSR_14 gnd vdd FILL
XFILL_61_DFFSR_9 gnd vdd FILL
XFILL_9_MUX2X1_114 gnd vdd FILL
XFILL_20_DFFSR_25 gnd vdd FILL
XFILL_20_DFFSR_36 gnd vdd FILL
XFILL_59_DFFSR_112 gnd vdd FILL
XFILL_9_MUX2X1_125 gnd vdd FILL
XFILL_59_DFFSR_123 gnd vdd FILL
XFILL_20_DFFSR_47 gnd vdd FILL
XFILL_59_DFFSR_134 gnd vdd FILL
XFILL_9_MUX2X1_136 gnd vdd FILL
XFILL_11_BUFX4_90 gnd vdd FILL
XFILL_20_DFFSR_58 gnd vdd FILL
XFILL_59_DFFSR_145 gnd vdd FILL
XFILL_9_MUX2X1_147 gnd vdd FILL
XFILL_59_DFFSR_156 gnd vdd FILL
XFILL_9_MUX2X1_158 gnd vdd FILL
XFILL_20_DFFSR_69 gnd vdd FILL
XFILL_9_MUX2X1_169 gnd vdd FILL
XFILL_59_DFFSR_167 gnd vdd FILL
XFILL_59_DFFSR_178 gnd vdd FILL
XFILL_60_DFFSR_13 gnd vdd FILL
XFILL_2_DFFSR_105 gnd vdd FILL
XFILL_6_OAI22X1_50 gnd vdd FILL
XFILL_59_DFFSR_189 gnd vdd FILL
XFILL_60_DFFSR_24 gnd vdd FILL
XFILL_2_DFFSR_116 gnd vdd FILL
XFILL_60_DFFSR_35 gnd vdd FILL
XFILL_2_DFFSR_127 gnd vdd FILL
XFILL_2_DFFSR_138 gnd vdd FILL
XFILL_60_DFFSR_46 gnd vdd FILL
XFILL_60_DFFSR_57 gnd vdd FILL
XFILL_2_DFFSR_149 gnd vdd FILL
XDFFSR_60 DFFSR_60/Q DFFSR_64/CLK DFFSR_69/R vdd DFFSR_60/D gnd vdd DFFSR
XFILL_60_DFFSR_68 gnd vdd FILL
XDFFSR_71 DFFSR_71/Q DFFSR_73/CLK DFFSR_73/R vdd DFFSR_71/D gnd vdd DFFSR
XDFFSR_82 DFFSR_82/Q DFFSR_84/CLK DFFSR_82/R vdd DFFSR_82/D gnd vdd DFFSR
XFILL_60_DFFSR_79 gnd vdd FILL
XDFFSR_93 DFFSR_93/Q DFFSR_93/CLK DFFSR_93/R vdd DFFSR_93/D gnd vdd DFFSR
XFILL_6_DFFSR_104 gnd vdd FILL
XFILL_10_MUX2X1_13 gnd vdd FILL
XFILL_6_DFFSR_115 gnd vdd FILL
XFILL_6_DFFSR_126 gnd vdd FILL
XFILL_3_DFFSR_15 gnd vdd FILL
XFILL_10_MUX2X1_24 gnd vdd FILL
XFILL_6_DFFSR_137 gnd vdd FILL
XFILL_10_MUX2X1_35 gnd vdd FILL
XFILL_3_DFFSR_26 gnd vdd FILL
XFILL_1_BUFX4_4 gnd vdd FILL
XFILL_6_DFFSR_148 gnd vdd FILL
XFILL_3_DFFSR_37 gnd vdd FILL
XFILL_10_MUX2X1_46 gnd vdd FILL
XFILL_3_DFFSR_48 gnd vdd FILL
XFILL_14_BUFX4_2 gnd vdd FILL
XFILL_6_DFFSR_159 gnd vdd FILL
XFILL_10_MUX2X1_57 gnd vdd FILL
XFILL_10_MUX2X1_68 gnd vdd FILL
XFILL_3_DFFSR_59 gnd vdd FILL
XFILL_10_MUX2X1_79 gnd vdd FILL
XFILL_6_3_0 gnd vdd FILL
XFILL_40_DFFSR_190 gnd vdd FILL
XFILL_14_MUX2X1_12 gnd vdd FILL
XFILL_14_MUX2X1_23 gnd vdd FILL
XFILL_5_INVX1_80 gnd vdd FILL
XFILL_14_MUX2X1_34 gnd vdd FILL
XFILL_5_INVX1_91 gnd vdd FILL
XFILL_14_MUX2X1_45 gnd vdd FILL
XFILL_14_MUX2X1_56 gnd vdd FILL
XFILL_14_MUX2X1_67 gnd vdd FILL
XFILL_2_NOR3X1_16 gnd vdd FILL
XFILL_14_MUX2X1_78 gnd vdd FILL
XFILL_12_MUX2X1_1 gnd vdd FILL
XFILL_14_MUX2X1_89 gnd vdd FILL
XFILL_2_NOR3X1_27 gnd vdd FILL
XFILL_18_MUX2X1_11 gnd vdd FILL
XFILL_2_NOR3X1_38 gnd vdd FILL
XFILL_18_MUX2X1_22 gnd vdd FILL
XFILL_2_NOR3X1_49 gnd vdd FILL
XFILL_18_MUX2X1_33 gnd vdd FILL
XFILL_18_MUX2X1_44 gnd vdd FILL
XFILL_18_MUX2X1_55 gnd vdd FILL
XFILL_0_INVX1_8 gnd vdd FILL
XFILL_18_MUX2X1_66 gnd vdd FILL
XFILL_15_7_1 gnd vdd FILL
XFILL_18_MUX2X1_77 gnd vdd FILL
XFILL_6_NOR3X1_15 gnd vdd FILL
XFILL_18_MUX2X1_88 gnd vdd FILL
XFILL_6_NOR3X1_26 gnd vdd FILL
XFILL_18_MUX2X1_99 gnd vdd FILL
XFILL_14_2_0 gnd vdd FILL
XFILL_6_NOR3X1_37 gnd vdd FILL
XFILL_22_DFFSR_102 gnd vdd FILL
XFILL_6_NOR3X1_48 gnd vdd FILL
XFILL_22_DFFSR_113 gnd vdd FILL
XFILL_22_DFFSR_124 gnd vdd FILL
XFILL_22_DFFSR_135 gnd vdd FILL
XFILL_22_DFFSR_146 gnd vdd FILL
XFILL_22_DFFSR_157 gnd vdd FILL
XFILL_22_DFFSR_168 gnd vdd FILL
XFILL_22_DFFSR_179 gnd vdd FILL
XFILL_26_DFFSR_101 gnd vdd FILL
XFILL_3_INVX1_108 gnd vdd FILL
XFILL_3_INVX1_119 gnd vdd FILL
XFILL_26_DFFSR_112 gnd vdd FILL
XFILL_1_NAND3X1_17 gnd vdd FILL
XFILL_26_DFFSR_123 gnd vdd FILL
XFILL_26_DFFSR_134 gnd vdd FILL
XFILL_1_NAND3X1_28 gnd vdd FILL
XFILL_26_DFFSR_145 gnd vdd FILL
XFILL_1_NAND3X1_39 gnd vdd FILL
XFILL_26_DFFSR_156 gnd vdd FILL
XINVX1_110 DFFSR_68/Q gnd NOR2X1_60/A vdd INVX1
XFILL_26_DFFSR_167 gnd vdd FILL
XFILL_5_NAND2X1_19 gnd vdd FILL
XFILL_26_DFFSR_178 gnd vdd FILL
XFILL_5_NOR2X1_2 gnd vdd FILL
XFILL_7_INVX1_107 gnd vdd FILL
XFILL_26_DFFSR_189 gnd vdd FILL
XINVX1_121 INVX1_121/A gnd INVX1_121/Y vdd INVX1
XFILL_7_INVX1_118 gnd vdd FILL
XINVX1_132 INVX1_132/A gnd INVX1_132/Y vdd INVX1
XFILL_7_INVX1_129 gnd vdd FILL
XINVX1_143 INVX1_143/A gnd OAI22X1_4/A vdd INVX1
XINVX1_154 INVX1_154/A gnd NOR2X1_98/A vdd INVX1
XINVX1_165 INVX1_165/A gnd OAI21X1_2/A vdd INVX1
XFILL_4_INVX8_2 gnd vdd FILL
XINVX1_176 INVX1_176/A gnd INVX1_176/Y vdd INVX1
XINVX1_187 INVX1_187/A gnd INVX1_187/Y vdd INVX1
XINVX1_198 DFFSR_91/Q gnd INVX1_198/Y vdd INVX1
XFILL_15_MUX2X1_150 gnd vdd FILL
XFILL_29_DFFSR_80 gnd vdd FILL
XFILL_22_NOR3X1_13 gnd vdd FILL
XFILL_15_MUX2X1_161 gnd vdd FILL
XFILL_22_NOR3X1_24 gnd vdd FILL
XFILL_29_DFFSR_91 gnd vdd FILL
XFILL_15_MUX2X1_172 gnd vdd FILL
XFILL_22_NOR3X1_35 gnd vdd FILL
XFILL_15_MUX2X1_183 gnd vdd FILL
XFILL_72_DFFSR_202 gnd vdd FILL
XFILL_22_NOR3X1_46 gnd vdd FILL
XFILL_15_MUX2X1_194 gnd vdd FILL
XFILL_72_DFFSR_213 gnd vdd FILL
XFILL_72_DFFSR_224 gnd vdd FILL
XFILL_72_DFFSR_235 gnd vdd FILL
XFILL_72_DFFSR_246 gnd vdd FILL
XFILL_26_NOR3X1_12 gnd vdd FILL
XFILL_21_DFFSR_2 gnd vdd FILL
XFILL_72_DFFSR_257 gnd vdd FILL
XFILL_72_DFFSR_268 gnd vdd FILL
XFILL_69_DFFSR_90 gnd vdd FILL
XFILL_26_NOR3X1_23 gnd vdd FILL
XFILL_26_NOR3X1_34 gnd vdd FILL
XFILL_65_6_1 gnd vdd FILL
XFILL_76_DFFSR_201 gnd vdd FILL
XFILL_26_NOR3X1_45 gnd vdd FILL
XFILL_76_DFFSR_212 gnd vdd FILL
XFILL_64_1_0 gnd vdd FILL
XFILL_76_DFFSR_223 gnd vdd FILL
XFILL_76_DFFSR_234 gnd vdd FILL
XFILL_1_NOR3X1_6 gnd vdd FILL
XFILL_76_DFFSR_245 gnd vdd FILL
XFILL_76_DFFSR_256 gnd vdd FILL
XFILL_76_DFFSR_267 gnd vdd FILL
XFILL_31_CLKBUF1_8 gnd vdd FILL
XFILL_34_1 gnd vdd FILL
XFILL_9_AOI21X1_19 gnd vdd FILL
XFILL_35_CLKBUF1_7 gnd vdd FILL
XFILL_20_CLKBUF1_18 gnd vdd FILL
XFILL_20_CLKBUF1_29 gnd vdd FILL
XFILL_43_DFFSR_6 gnd vdd FILL
XFILL_1_NOR2X1_107 gnd vdd FILL
XFILL_1_NOR2X1_118 gnd vdd FILL
XFILL_1_NOR2X1_129 gnd vdd FILL
XFILL_11_NAND2X1_11 gnd vdd FILL
XFILL_8_BUFX4_19 gnd vdd FILL
XFILL_11_NAND2X1_22 gnd vdd FILL
XFILL_11_NAND2X1_33 gnd vdd FILL
XFILL_11_NAND2X1_44 gnd vdd FILL
XFILL_11_NAND2X1_55 gnd vdd FILL
XFILL_1_OAI21X1_3 gnd vdd FILL
XFILL_56_6_1 gnd vdd FILL
XFILL_11_NAND2X1_66 gnd vdd FILL
XFILL_9_OAI22X1_16 gnd vdd FILL
XFILL_11_NAND2X1_77 gnd vdd FILL
XFILL_11_NAND2X1_88 gnd vdd FILL
XFILL_9_OAI22X1_27 gnd vdd FILL
XFILL_55_1_0 gnd vdd FILL
XFILL_9_OAI22X1_38 gnd vdd FILL
XFILL_9_OAI22X1_49 gnd vdd FILL
XFILL_43_DFFSR_201 gnd vdd FILL
XFILL_43_DFFSR_212 gnd vdd FILL
XFILL_5_OAI21X1_2 gnd vdd FILL
XFILL_43_DFFSR_223 gnd vdd FILL
XFILL_43_DFFSR_234 gnd vdd FILL
XFILL_2_NOR2X1_60 gnd vdd FILL
XFILL_43_DFFSR_245 gnd vdd FILL
XFILL_43_DFFSR_256 gnd vdd FILL
XFILL_43_DFFSR_267 gnd vdd FILL
XFILL_2_NOR2X1_71 gnd vdd FILL
XNAND3X1_107 NOR2X1_5/A BUFX4_7/Y AND2X2_4/A gnd OAI21X1_18/C vdd NAND3X1
XFILL_8_NAND3X1_70 gnd vdd FILL
XFILL_2_NOR2X1_82 gnd vdd FILL
XFILL_2_NOR2X1_93 gnd vdd FILL
XNAND3X1_118 NAND3X1_118/A NAND3X1_118/B NAND3X1_118/C gnd NOR3X1_31/C vdd NAND3X1
XFILL_8_NAND3X1_81 gnd vdd FILL
XFILL_70_DFFSR_101 gnd vdd FILL
XFILL_8_NAND3X1_92 gnd vdd FILL
XFILL_47_DFFSR_200 gnd vdd FILL
XNAND3X1_129 DFFSR_141/Q BUFX4_92/Y AND2X2_4/A gnd OAI21X1_21/C vdd NAND3X1
XFILL_47_DFFSR_211 gnd vdd FILL
XFILL_70_DFFSR_112 gnd vdd FILL
XFILL_5_BUFX4_5 gnd vdd FILL
XFILL_47_DFFSR_222 gnd vdd FILL
XFILL_9_OAI21X1_1 gnd vdd FILL
XFILL_70_DFFSR_123 gnd vdd FILL
XFILL_70_DFFSR_134 gnd vdd FILL
XFILL_47_DFFSR_233 gnd vdd FILL
XFILL_70_DFFSR_145 gnd vdd FILL
XFILL_47_DFFSR_244 gnd vdd FILL
XFILL_70_DFFSR_156 gnd vdd FILL
XFILL_47_DFFSR_255 gnd vdd FILL
XFILL_6_NOR2X1_70 gnd vdd FILL
XFILL_70_DFFSR_167 gnd vdd FILL
XFILL_15_AND2X2_7 gnd vdd FILL
XFILL_47_DFFSR_266 gnd vdd FILL
XFILL_70_DFFSR_178 gnd vdd FILL
XFILL_6_NOR2X1_81 gnd vdd FILL
XFILL_6_NOR2X1_92 gnd vdd FILL
XFILL_2_OAI21X1_18 gnd vdd FILL
XFILL_74_DFFSR_100 gnd vdd FILL
XFILL_70_DFFSR_189 gnd vdd FILL
XFILL_2_OAI21X1_29 gnd vdd FILL
XFILL_74_DFFSR_111 gnd vdd FILL
XFILL_74_DFFSR_122 gnd vdd FILL
XFILL_74_DFFSR_133 gnd vdd FILL
XFILL_74_DFFSR_144 gnd vdd FILL
XFILL_15_AOI21X1_11 gnd vdd FILL
XFILL_74_DFFSR_155 gnd vdd FILL
XFILL_15_AOI21X1_22 gnd vdd FILL
XFILL_15_AOI21X1_33 gnd vdd FILL
XFILL_74_DFFSR_166 gnd vdd FILL
XFILL_15_AOI21X1_44 gnd vdd FILL
XFILL_74_DFFSR_177 gnd vdd FILL
XFILL_74_DFFSR_188 gnd vdd FILL
XFILL_15_AOI21X1_55 gnd vdd FILL
XFILL_1_NAND2X1_50 gnd vdd FILL
XFILL_78_DFFSR_110 gnd vdd FILL
XFILL_74_DFFSR_199 gnd vdd FILL
XFILL_12_BUFX4_13 gnd vdd FILL
XFILL_15_AOI21X1_66 gnd vdd FILL
XFILL_1_NAND2X1_61 gnd vdd FILL
XFILL_1_NAND2X1_72 gnd vdd FILL
XFILL_15_AOI21X1_77 gnd vdd FILL
XFILL_78_DFFSR_121 gnd vdd FILL
XFILL_78_DFFSR_132 gnd vdd FILL
XFILL_12_BUFX4_24 gnd vdd FILL
XFILL_4_INVX1_9 gnd vdd FILL
XFILL_78_DFFSR_143 gnd vdd FILL
XFILL_12_BUFX4_35 gnd vdd FILL
XFILL_1_NAND2X1_83 gnd vdd FILL
XFILL_78_DFFSR_154 gnd vdd FILL
XFILL_12_BUFX4_46 gnd vdd FILL
XFILL_1_NAND2X1_94 gnd vdd FILL
XFILL_12_BUFX4_57 gnd vdd FILL
XFILL_78_DFFSR_165 gnd vdd FILL
XFILL_12_BUFX4_68 gnd vdd FILL
XFILL_78_DFFSR_176 gnd vdd FILL
XFILL_1_BUFX2_1 gnd vdd FILL
XFILL_78_DFFSR_187 gnd vdd FILL
XFILL_12_BUFX4_79 gnd vdd FILL
XFILL_78_DFFSR_198 gnd vdd FILL
XFILL_2_NAND2X1_4 gnd vdd FILL
XFILL_47_6_1 gnd vdd FILL
XFILL_46_1_0 gnd vdd FILL
XFILL_6_NAND2X1_3 gnd vdd FILL
XFILL_6_INVX1_14 gnd vdd FILL
XFILL_10_DFFSR_201 gnd vdd FILL
XFILL_6_INVX1_25 gnd vdd FILL
XFILL_6_INVX1_36 gnd vdd FILL
XFILL_10_DFFSR_212 gnd vdd FILL
XFILL_18_MUX2X1_105 gnd vdd FILL
XFILL_8_INVX8_3 gnd vdd FILL
XFILL_6_INVX1_47 gnd vdd FILL
XFILL_18_MUX2X1_116 gnd vdd FILL
XFILL_10_DFFSR_223 gnd vdd FILL
XFILL_7_AND2X2_6 gnd vdd FILL
XFILL_10_DFFSR_234 gnd vdd FILL
XFILL_18_MUX2X1_127 gnd vdd FILL
XFILL_6_INVX1_58 gnd vdd FILL
XFILL_18_MUX2X1_138 gnd vdd FILL
XFILL_6_INVX1_69 gnd vdd FILL
XFILL_10_DFFSR_245 gnd vdd FILL
XFILL_18_MUX2X1_149 gnd vdd FILL
XFILL_5_AOI21X1_50 gnd vdd FILL
XFILL_10_DFFSR_256 gnd vdd FILL
XFILL_5_AOI21X1_61 gnd vdd FILL
XFILL_10_DFFSR_267 gnd vdd FILL
XFILL_5_AOI21X1_72 gnd vdd FILL
XFILL_15_OAI22X1_30 gnd vdd FILL
XFILL_15_OAI22X1_41 gnd vdd FILL
XFILL_14_DFFSR_200 gnd vdd FILL
XFILL_30_5_1 gnd vdd FILL
XFILL_14_DFFSR_211 gnd vdd FILL
XFILL_14_DFFSR_222 gnd vdd FILL
XFILL_14_DFFSR_233 gnd vdd FILL
XFILL_14_DFFSR_244 gnd vdd FILL
XFILL_25_DFFSR_3 gnd vdd FILL
XDFFSR_105 NAND3X1_3/A DFFSR_78/CLK DFFSR_78/R vdd DFFSR_105/D gnd vdd DFFSR
XFILL_14_DFFSR_255 gnd vdd FILL
XFILL_4_BUFX4_12 gnd vdd FILL
XFILL_8_NOR2X1_160 gnd vdd FILL
XDFFSR_116 INVX1_187/A CLKBUF1_31/Y DFFSR_64/R vdd DFFSR_116/D gnd vdd DFFSR
XFILL_14_DFFSR_266 gnd vdd FILL
XFILL_82_DFFSR_4 gnd vdd FILL
XFILL_4_BUFX4_23 gnd vdd FILL
XFILL_41_DFFSR_100 gnd vdd FILL
XDFFSR_127 INVX1_171/A DFFSR_64/CLK DFFSR_2/R vdd DFFSR_127/D gnd vdd DFFSR
XFILL_8_NOR2X1_171 gnd vdd FILL
XFILL_4_BUFX4_34 gnd vdd FILL
XDFFSR_138 INVX1_164/A DFFSR_55/CLK DFFSR_55/R vdd DFFSR_138/D gnd vdd DFFSR
XFILL_8_NOR2X1_182 gnd vdd FILL
XFILL_4_BUFX4_45 gnd vdd FILL
XDFFSR_149 DFFSR_149/Q CLKBUF1_6/Y DFFSR_48/R vdd DFFSR_149/D gnd vdd DFFSR
XFILL_18_DFFSR_210 gnd vdd FILL
XFILL_8_NOR2X1_193 gnd vdd FILL
XFILL_41_DFFSR_111 gnd vdd FILL
XFILL_18_DFFSR_221 gnd vdd FILL
XFILL_4_BUFX4_56 gnd vdd FILL
XFILL_41_DFFSR_122 gnd vdd FILL
XFILL_1_INVX2_1 gnd vdd FILL
XFILL_2_AOI21X1_9 gnd vdd FILL
XFILL_41_DFFSR_133 gnd vdd FILL
XFILL_4_BUFX4_67 gnd vdd FILL
XFILL_41_DFFSR_144 gnd vdd FILL
XFILL_4_BUFX4_78 gnd vdd FILL
XFILL_18_DFFSR_232 gnd vdd FILL
XFILL_18_DFFSR_243 gnd vdd FILL
XFILL_4_BUFX4_89 gnd vdd FILL
XFILL_41_DFFSR_155 gnd vdd FILL
XFILL_18_DFFSR_254 gnd vdd FILL
XFILL_41_DFFSR_166 gnd vdd FILL
XFILL_18_DFFSR_265 gnd vdd FILL
XFILL_41_DFFSR_177 gnd vdd FILL
XFILL_41_DFFSR_188 gnd vdd FILL
XFILL_41_DFFSR_199 gnd vdd FILL
XFILL_45_DFFSR_110 gnd vdd FILL
XFILL_45_DFFSR_121 gnd vdd FILL
XFILL_45_DFFSR_132 gnd vdd FILL
XFILL_6_AOI21X1_8 gnd vdd FILL
XFILL_45_DFFSR_143 gnd vdd FILL
XFILL_45_DFFSR_154 gnd vdd FILL
XFILL_45_DFFSR_165 gnd vdd FILL
XFILL_45_DFFSR_176 gnd vdd FILL
XFILL_8_MUX2X1_100 gnd vdd FILL
XFILL_45_DFFSR_187 gnd vdd FILL
XFILL_8_MUX2X1_111 gnd vdd FILL
XFILL_45_DFFSR_198 gnd vdd FILL
XFILL_8_MUX2X1_122 gnd vdd FILL
XFILL_49_DFFSR_120 gnd vdd FILL
XFILL_49_DFFSR_131 gnd vdd FILL
XFILL_47_DFFSR_7 gnd vdd FILL
XFILL_8_MUX2X1_133 gnd vdd FILL
XFILL_8_MUX2X1_144 gnd vdd FILL
XFILL_49_DFFSR_142 gnd vdd FILL
XNOR3X1_16 INVX1_79/Y NOR3X1_49/B NOR3X1_39/C gnd NOR3X1_17/C vdd NOR3X1
XFILL_8_MUX2X1_155 gnd vdd FILL
XFILL_49_DFFSR_153 gnd vdd FILL
XFILL_11_AOI22X1_5 gnd vdd FILL
XNOR3X1_27 NOR3X1_27/A NOR3X1_27/B NOR3X1_27/C gnd NOR3X1_27/Y vdd NOR3X1
XFILL_38_6_1 gnd vdd FILL
XFILL_8_MUX2X1_166 gnd vdd FILL
XFILL_49_DFFSR_164 gnd vdd FILL
XNOR3X1_38 NOR3X1_38/A NOR3X1_38/B NOR3X1_38/C gnd NOR3X1_38/Y vdd NOR3X1
XFILL_8_MUX2X1_177 gnd vdd FILL
XNOR3X1_49 NOR3X1_49/A NOR3X1_49/B NOR3X1_6/B gnd NOR3X1_50/C vdd NOR3X1
XFILL_49_DFFSR_175 gnd vdd FILL
XFILL_37_1_0 gnd vdd FILL
XFILL_49_DFFSR_186 gnd vdd FILL
XFILL_8_MUX2X1_188 gnd vdd FILL
XFILL_49_DFFSR_197 gnd vdd FILL
XFILL_15_AOI22X1_4 gnd vdd FILL
XFILL_10_NAND3X1_19 gnd vdd FILL
XFILL_19_AOI22X1_3 gnd vdd FILL
XFILL_21_5_1 gnd vdd FILL
XFILL_20_0_0 gnd vdd FILL
XFILL_39_DFFSR_12 gnd vdd FILL
XFILL_30_CLKBUF1_19 gnd vdd FILL
XFILL_39_DFFSR_23 gnd vdd FILL
XFILL_39_DFFSR_34 gnd vdd FILL
XFILL_39_DFFSR_45 gnd vdd FILL
XFILL_39_DFFSR_56 gnd vdd FILL
XFILL_39_DFFSR_67 gnd vdd FILL
XFILL_39_DFFSR_78 gnd vdd FILL
XFILL_39_DFFSR_89 gnd vdd FILL
XFILL_79_DFFSR_11 gnd vdd FILL
XFILL_79_DFFSR_22 gnd vdd FILL
XFILL_79_DFFSR_33 gnd vdd FILL
XFILL_79_DFFSR_44 gnd vdd FILL
XFILL_0_DFFSR_19 gnd vdd FILL
XFILL_79_DFFSR_55 gnd vdd FILL
XFILL_79_DFFSR_66 gnd vdd FILL
XFILL_79_DFFSR_77 gnd vdd FILL
XFILL_10_NOR2X1_7 gnd vdd FILL
XFILL_79_DFFSR_88 gnd vdd FILL
XFILL_79_DFFSR_99 gnd vdd FILL
XFILL_2_INVX1_40 gnd vdd FILL
XFILL_12_DFFSR_110 gnd vdd FILL
XFILL_2_INVX1_51 gnd vdd FILL
XFILL_9_BUFX4_6 gnd vdd FILL
XFILL_2_INVX1_62 gnd vdd FILL
XFILL_12_DFFSR_121 gnd vdd FILL
XFILL_12_DFFSR_132 gnd vdd FILL
XFILL_12_DFFSR_143 gnd vdd FILL
XFILL_48_DFFSR_10 gnd vdd FILL
XFILL_2_INVX1_73 gnd vdd FILL
XFILL_12_DFFSR_154 gnd vdd FILL
XFILL_48_DFFSR_21 gnd vdd FILL
XFILL_2_INVX1_84 gnd vdd FILL
XFILL_2_INVX1_95 gnd vdd FILL
XFILL_48_DFFSR_32 gnd vdd FILL
XFILL_12_DFFSR_165 gnd vdd FILL
XFILL_19_NOR3X1_7 gnd vdd FILL
XFILL_48_DFFSR_43 gnd vdd FILL
XFILL_1_CLKBUF1_8 gnd vdd FILL
XFILL_12_DFFSR_176 gnd vdd FILL
XFILL_12_DFFSR_187 gnd vdd FILL
XFILL_48_DFFSR_54 gnd vdd FILL
XFILL_12_DFFSR_198 gnd vdd FILL
XFILL_48_DFFSR_65 gnd vdd FILL
XFILL_48_DFFSR_76 gnd vdd FILL
XFILL_29_6_1 gnd vdd FILL
XFILL_16_DFFSR_120 gnd vdd FILL
XFILL_0_NAND3X1_14 gnd vdd FILL
XFILL_48_DFFSR_87 gnd vdd FILL
XFILL_4_6_1 gnd vdd FILL
XFILL_16_DFFSR_131 gnd vdd FILL
XFILL_0_NAND3X1_25 gnd vdd FILL
XFILL_48_DFFSR_98 gnd vdd FILL
XFILL_16_DFFSR_142 gnd vdd FILL
XFILL_0_NAND3X1_36 gnd vdd FILL
XFILL_28_1_0 gnd vdd FILL
XFILL_16_DFFSR_153 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XFILL_0_NAND3X1_47 gnd vdd FILL
XFILL_0_NAND3X1_58 gnd vdd FILL
XFILL_4_NAND2X1_16 gnd vdd FILL
XFILL_16_DFFSR_164 gnd vdd FILL
XFILL_5_CLKBUF1_7 gnd vdd FILL
XFILL_0_NAND3X1_69 gnd vdd FILL
XFILL_16_DFFSR_175 gnd vdd FILL
XFILL_4_NAND2X1_27 gnd vdd FILL
XFILL_16_DFFSR_186 gnd vdd FILL
XFILL_16_DFFSR_197 gnd vdd FILL
XFILL_17_DFFSR_20 gnd vdd FILL
XFILL_4_NAND2X1_38 gnd vdd FILL
XFILL_4_NAND2X1_49 gnd vdd FILL
XFILL_0_BUFX4_60 gnd vdd FILL
XFILL_17_DFFSR_31 gnd vdd FILL
XFILL_0_BUFX4_71 gnd vdd FILL
XFILL_17_DFFSR_42 gnd vdd FILL
XFILL_0_BUFX4_82 gnd vdd FILL
XFILL_0_BUFX4_93 gnd vdd FILL
XFILL_17_DFFSR_53 gnd vdd FILL
XFILL_1_BUFX4_102 gnd vdd FILL
XFILL_17_DFFSR_64 gnd vdd FILL
XFILL_17_DFFSR_75 gnd vdd FILL
XFILL_17_DFFSR_86 gnd vdd FILL
XFILL_12_NOR3X1_10 gnd vdd FILL
XFILL_17_DFFSR_97 gnd vdd FILL
XFILL_9_CLKBUF1_6 gnd vdd FILL
XFILL_12_NOR3X1_21 gnd vdd FILL
XFILL_5_BUFX2_2 gnd vdd FILL
XFILL_12_NOR3X1_32 gnd vdd FILL
XFILL_57_DFFSR_30 gnd vdd FILL
XFILL_14_MUX2X1_180 gnd vdd FILL
XFILL_57_DFFSR_41 gnd vdd FILL
XFILL_12_5_1 gnd vdd FILL
XFILL_12_NOR3X1_43 gnd vdd FILL
XFILL_28_NOR3X1_5 gnd vdd FILL
XFILL_14_MUX2X1_191 gnd vdd FILL
XFILL_62_DFFSR_210 gnd vdd FILL
XFILL_57_DFFSR_52 gnd vdd FILL
XFILL_62_DFFSR_221 gnd vdd FILL
XFILL_57_DFFSR_63 gnd vdd FILL
XFILL_5_BUFX4_101 gnd vdd FILL
XFILL_11_0_0 gnd vdd FILL
XFILL_57_DFFSR_74 gnd vdd FILL
XFILL_62_DFFSR_232 gnd vdd FILL
XFILL_62_DFFSR_243 gnd vdd FILL
XFILL_57_DFFSR_85 gnd vdd FILL
XFILL_62_DFFSR_254 gnd vdd FILL
XFILL_57_DFFSR_96 gnd vdd FILL
XFILL_62_DFFSR_265 gnd vdd FILL
XFILL_16_NOR3X1_20 gnd vdd FILL
XFILL_16_NOR3X1_31 gnd vdd FILL
XFILL_2_NOR2X1_6 gnd vdd FILL
XFILL_16_NOR3X1_42 gnd vdd FILL
XFILL_64_DFFSR_1 gnd vdd FILL
XFILL_66_DFFSR_220 gnd vdd FILL
XFILL_10_NOR2X1_109 gnd vdd FILL
XFILL_66_DFFSR_231 gnd vdd FILL
XFILL_9_BUFX4_100 gnd vdd FILL
XFILL_26_DFFSR_40 gnd vdd FILL
XFILL_66_DFFSR_242 gnd vdd FILL
XFILL_26_DFFSR_51 gnd vdd FILL
XFILL_66_DFFSR_253 gnd vdd FILL
XFILL_26_DFFSR_62 gnd vdd FILL
XFILL_66_DFFSR_264 gnd vdd FILL
XFILL_66_DFFSR_275 gnd vdd FILL
XFILL_21_CLKBUF1_5 gnd vdd FILL
XFILL_26_DFFSR_73 gnd vdd FILL
XFILL_26_DFFSR_84 gnd vdd FILL
XFILL_26_DFFSR_95 gnd vdd FILL
XFILL_8_AOI21X1_16 gnd vdd FILL
XFILL_8_AOI21X1_27 gnd vdd FILL
XFILL_1_MUX2X1_4 gnd vdd FILL
XFILL_8_AOI21X1_38 gnd vdd FILL
XFILL_8_AOI21X1_49 gnd vdd FILL
XFILL_66_DFFSR_50 gnd vdd FILL
XFILL_66_DFFSR_61 gnd vdd FILL
XFILL_18_OAI22X1_18 gnd vdd FILL
XFILL_25_CLKBUF1_4 gnd vdd FILL
XFILL_66_DFFSR_72 gnd vdd FILL
XFILL_18_OAI22X1_29 gnd vdd FILL
XFILL_66_DFFSR_83 gnd vdd FILL
XFILL_3_NOR2X1_14 gnd vdd FILL
XFILL_66_DFFSR_94 gnd vdd FILL
XFILL_3_NOR2X1_25 gnd vdd FILL
XFILL_3_NOR2X1_36 gnd vdd FILL
XFILL_3_NOR2X1_47 gnd vdd FILL
XFILL_29_DFFSR_4 gnd vdd FILL
XNAND3X1_60 AND2X2_5/B AND2X2_6/A BUFX4_57/Y gnd NOR2X1_60/B vdd NAND3X1
XFILL_3_NOR2X1_58 gnd vdd FILL
XNAND3X1_71 NOR2X1_79/A BUFX4_88/Y NOR2X1_36/Y gnd OAI21X1_4/C vdd NAND3X1
XFILL_9_DFFSR_30 gnd vdd FILL
XFILL_86_DFFSR_5 gnd vdd FILL
XFILL_2_CLKBUF1_19 gnd vdd FILL
XFILL_3_NOR2X1_69 gnd vdd FILL
XNAND3X1_82 NAND3X1_82/A NAND3X1_82/B NAND3X1_82/C gnd NOR2X1_61/B vdd NAND3X1
XFILL_9_DFFSR_41 gnd vdd FILL
XFILL_29_CLKBUF1_3 gnd vdd FILL
XNAND3X1_93 NOR2X1_90/A BUFX4_88/Y NOR2X1_36/Y gnd OAI21X1_14/C vdd NAND3X1
XFILL_9_DFFSR_52 gnd vdd FILL
XFILL_9_DFFSR_63 gnd vdd FILL
XFILL_19_1_0 gnd vdd FILL
XFILL_7_NAND3X1_130 gnd vdd FILL
XFILL_7_NOR2X1_13 gnd vdd FILL
XFILL_5_INVX2_2 gnd vdd FILL
XFILL_9_DFFSR_74 gnd vdd FILL
XFILL_48_DFFSR_209 gnd vdd FILL
XFILL_9_DFFSR_85 gnd vdd FILL
XFILL_35_DFFSR_60 gnd vdd FILL
XFILL_7_NOR2X1_24 gnd vdd FILL
XFILL_9_DFFSR_96 gnd vdd FILL
XFILL_7_NOR2X1_35 gnd vdd FILL
XFILL_35_DFFSR_71 gnd vdd FILL
XFILL_35_DFFSR_82 gnd vdd FILL
XNOR2X1_60 NOR2X1_60/A NOR2X1_60/B gnd NOR3X1_13/A vdd NOR2X1
XFILL_7_NOR2X1_46 gnd vdd FILL
XFILL_11_OAI22X1_8 gnd vdd FILL
XNOR2X1_71 INVX1_77/Y OAI22X1_1/D gnd NOR3X1_25/A vdd NOR2X1
XFILL_7_NOR2X1_57 gnd vdd FILL
XFILL_62_4_1 gnd vdd FILL
XFILL_35_DFFSR_93 gnd vdd FILL
XFILL_7_NOR2X1_68 gnd vdd FILL
XNOR2X1_82 NOR2X1_82/A NOR2X1_82/B gnd NOR2X1_82/Y vdd NOR2X1
XFILL_7_NOR2X1_79 gnd vdd FILL
XNOR2X1_93 NOR2X1_93/A NOR2X1_93/B gnd NOR2X1_93/Y vdd NOR2X1
XFILL_0_NOR2X1_104 gnd vdd FILL
XFILL_75_DFFSR_109 gnd vdd FILL
XFILL_0_NOR2X1_115 gnd vdd FILL
XFILL_0_NOR2X1_126 gnd vdd FILL
XFILL_75_DFFSR_70 gnd vdd FILL
XFILL_75_DFFSR_81 gnd vdd FILL
XFILL_0_NOR2X1_137 gnd vdd FILL
XFILL_75_DFFSR_92 gnd vdd FILL
XFILL_15_OAI22X1_7 gnd vdd FILL
XFILL_0_NOR2X1_148 gnd vdd FILL
XFILL_0_NOR2X1_159 gnd vdd FILL
XFILL_11_3 gnd vdd FILL
XFILL_79_DFFSR_108 gnd vdd FILL
XFILL_10_NAND2X1_30 gnd vdd FILL
XFILL_10_NAND2X1_41 gnd vdd FILL
XFILL_79_DFFSR_119 gnd vdd FILL
XFILL_10_NAND2X1_52 gnd vdd FILL
XFILL_19_OAI22X1_6 gnd vdd FILL
XFILL_10_NAND2X1_63 gnd vdd FILL
XFILL_8_OAI22X1_13 gnd vdd FILL
XFILL_10_NAND2X1_74 gnd vdd FILL
XFILL_8_OAI22X1_24 gnd vdd FILL
XFILL_10_NAND2X1_85 gnd vdd FILL
XFILL_8_OAI22X1_35 gnd vdd FILL
XFILL_10_NAND2X1_96 gnd vdd FILL
XFILL_44_DFFSR_80 gnd vdd FILL
XFILL_8_OAI22X1_46 gnd vdd FILL
XFILL_44_DFFSR_91 gnd vdd FILL
XBUFX2_9 BUFX2_9/A gnd addr[5] vdd BUFX2
XFILL_33_DFFSR_220 gnd vdd FILL
XFILL_33_DFFSR_231 gnd vdd FILL
XFILL_33_DFFSR_242 gnd vdd FILL
XFILL_33_DFFSR_253 gnd vdd FILL
XFILL_33_DFFSR_264 gnd vdd FILL
XFILL_33_DFFSR_275 gnd vdd FILL
XFILL_84_DFFSR_90 gnd vdd FILL
XFILL_5_NOR2X1_204 gnd vdd FILL
XFILL_60_DFFSR_120 gnd vdd FILL
XFILL_60_DFFSR_131 gnd vdd FILL
XFILL_37_DFFSR_230 gnd vdd FILL
XFILL_13_DFFSR_90 gnd vdd FILL
XFILL_60_DFFSR_142 gnd vdd FILL
XFILL_60_DFFSR_153 gnd vdd FILL
XFILL_37_DFFSR_241 gnd vdd FILL
XFILL_37_DFFSR_252 gnd vdd FILL
XFILL_3_MUX2X1_10 gnd vdd FILL
XNAND2X1_4 OAI21X1_1/A NAND2X1_4/B gnd NOR2X1_7/B vdd NAND2X1
XFILL_37_DFFSR_263 gnd vdd FILL
XFILL_60_DFFSR_164 gnd vdd FILL
XFILL_37_DFFSR_274 gnd vdd FILL
XFILL_60_DFFSR_175 gnd vdd FILL
XFILL_3_MUX2X1_21 gnd vdd FILL
XFILL_1_OAI21X1_15 gnd vdd FILL
XFILL_60_DFFSR_186 gnd vdd FILL
XFILL_19_CLKBUF1_11 gnd vdd FILL
XFILL_1_OAI21X1_26 gnd vdd FILL
XFILL_60_DFFSR_197 gnd vdd FILL
XFILL_3_MUX2X1_32 gnd vdd FILL
XFILL_1_OAI21X1_37 gnd vdd FILL
XFILL_3_MUX2X1_43 gnd vdd FILL
XFILL_19_CLKBUF1_22 gnd vdd FILL
XFILL_3_MUX2X1_54 gnd vdd FILL
XFILL_1_OAI21X1_48 gnd vdd FILL
XFILL_64_DFFSR_130 gnd vdd FILL
XFILL_19_CLKBUF1_33 gnd vdd FILL
XFILL_3_MUX2X1_65 gnd vdd FILL
XFILL_64_DFFSR_141 gnd vdd FILL
XFILL_64_DFFSR_152 gnd vdd FILL
XFILL_3_MUX2X1_76 gnd vdd FILL
XFILL_3_MUX2X1_87 gnd vdd FILL
XFILL_64_DFFSR_163 gnd vdd FILL
XFILL_14_AOI21X1_30 gnd vdd FILL
XFILL_3_MUX2X1_98 gnd vdd FILL
XFILL_64_DFFSR_174 gnd vdd FILL
XFILL_14_AOI21X1_41 gnd vdd FILL
XFILL_7_MUX2X1_20 gnd vdd FILL
XFILL_14_AOI21X1_52 gnd vdd FILL
XFILL_64_DFFSR_185 gnd vdd FILL
XFILL_7_MUX2X1_31 gnd vdd FILL
XFILL_14_AOI21X1_63 gnd vdd FILL
XFILL_64_DFFSR_196 gnd vdd FILL
XFILL_53_4_1 gnd vdd FILL
XFILL_7_MUX2X1_42 gnd vdd FILL
XFILL_15_DFFSR_209 gnd vdd FILL
XFILL_14_AOI21X1_74 gnd vdd FILL
XFILL_7_MUX2X1_53 gnd vdd FILL
XFILL_12_NAND3X1_9 gnd vdd FILL
XFILL_7_MUX2X1_64 gnd vdd FILL
XFILL_0_NAND2X1_80 gnd vdd FILL
XFILL_68_DFFSR_140 gnd vdd FILL
XNOR2X1_150 DFFSR_99/Q NOR2X1_153/B gnd NOR2X1_150/Y vdd NOR2X1
XNOR2X1_161 DFFSR_84/Q NOR2X1_161/B gnd NOR2X1_161/Y vdd NOR2X1
XFILL_7_MUX2X1_75 gnd vdd FILL
XFILL_68_DFFSR_151 gnd vdd FILL
XFILL_0_NAND2X1_91 gnd vdd FILL
XFILL_68_DFFSR_162 gnd vdd FILL
XFILL_7_MUX2X1_86 gnd vdd FILL
XFILL_7_MUX2X1_97 gnd vdd FILL
XFILL_68_DFFSR_173 gnd vdd FILL
XNOR2X1_172 NOR2X1_7/B INVX1_174/Y gnd MUX2X1_9/S vdd NOR2X1
XNOR2X1_183 DFFSR_25/Q MUX2X1_16/S gnd NOR2X1_183/Y vdd NOR2X1
XFILL_68_DFFSR_184 gnd vdd FILL
XNOR2X1_194 DFFSR_17/Q NOR2X1_195/B gnd NOR2X1_194/Y vdd NOR2X1
XFILL_68_DFFSR_195 gnd vdd FILL
XFILL_42_DFFSR_109 gnd vdd FILL
XFILL_19_DFFSR_208 gnd vdd FILL
XFILL_19_DFFSR_219 gnd vdd FILL
XFILL_46_DFFSR_108 gnd vdd FILL
XAOI21X1_9 BUFX4_67/Y AOI21X1_9/B AOI21X1_9/C gnd DFFSR_104/D vdd AOI21X1
XFILL_46_DFFSR_119 gnd vdd FILL
XMUX2X1_101 BUFX4_78/Y INVX1_148/Y NOR2X1_57/Y gnd DFFSR_163/D vdd MUX2X1
XMUX2X1_112 NOR2X1_98/A BUFX4_93/Y NAND2X1_23/Y gnd DFFSR_155/D vdd MUX2X1
XMUX2X1_123 BUFX4_68/Y INVX1_167/Y NOR2X1_136/Y gnd DFFSR_131/D vdd MUX2X1
XMUX2X1_134 INVX1_178/Y MUX2X1_7/B NAND2X1_2/Y gnd DFFSR_125/D vdd MUX2X1
XMUX2X1_145 BUFX4_67/Y INVX1_189/Y NOR2X1_142/Y gnd DFFSR_108/D vdd MUX2X1
XFILL_17_MUX2X1_102 gnd vdd FILL
XFILL_17_MUX2X1_113 gnd vdd FILL
XMUX2X1_156 BUFX4_99/Y INVX1_200/Y NOR2X1_155/Y gnd DFFSR_93/D vdd MUX2X1
XFILL_23_MUX2X1_40 gnd vdd FILL
XFILL_23_MUX2X1_51 gnd vdd FILL
XMUX2X1_167 BUFX4_67/Y INVX1_212/Y NOR2X1_164/Y gnd DFFSR_73/D vdd MUX2X1
XFILL_17_MUX2X1_124 gnd vdd FILL
XFILL_23_MUX2X1_62 gnd vdd FILL
XFILL_17_MUX2X1_135 gnd vdd FILL
XMUX2X1_178 BUFX4_93/Y INVX1_223/Y NOR2X1_166/Y gnd DFFSR_66/D vdd MUX2X1
XFILL_23_MUX2X1_73 gnd vdd FILL
XFILL_17_MUX2X1_146 gnd vdd FILL
XMUX2X1_189 BUFX4_67/Y INVX1_9/Y NOR2X1_169/Y gnd DFFSR_51/D vdd MUX2X1
XFILL_23_MUX2X1_84 gnd vdd FILL
XFILL_17_MUX2X1_157 gnd vdd FILL
XFILL_9_BUFX2_3 gnd vdd FILL
XFILL_23_MUX2X1_95 gnd vdd FILL
XFILL_17_MUX2X1_168 gnd vdd FILL
XFILL_4_AOI21X1_80 gnd vdd FILL
XFILL_17_MUX2X1_179 gnd vdd FILL
XINVX1_30 INVX1_30/A gnd INVX1_30/Y vdd INVX1
XINVX1_41 INVX1_41/A gnd INVX1_41/Y vdd INVX1
XFILL_30_DFFSR_4 gnd vdd FILL
XINVX1_52 INVX1_52/A gnd INVX1_52/Y vdd INVX1
XINVX1_63 INVX1_63/A gnd INVX1_63/Y vdd INVX1
XINVX1_74 INVX1_74/A gnd INVX1_74/Y vdd INVX1
XINVX1_85 INVX1_85/A gnd INVX1_85/Y vdd INVX1
XINVX1_96 INVX1_96/A gnd INVX1_96/Y vdd INVX1
XFILL_7_NOR2X1_190 gnd vdd FILL
XFILL_68_DFFSR_2 gnd vdd FILL
XFILL_31_DFFSR_130 gnd vdd FILL
XFILL_3_INVX1_18 gnd vdd FILL
XFILL_3_INVX1_29 gnd vdd FILL
XFILL_31_DFFSR_141 gnd vdd FILL
XFILL_31_DFFSR_152 gnd vdd FILL
XFILL_44_4_1 gnd vdd FILL
XFILL_31_DFFSR_163 gnd vdd FILL
XFILL_31_DFFSR_174 gnd vdd FILL
XFILL_31_DFFSR_185 gnd vdd FILL
XFILL_31_DFFSR_196 gnd vdd FILL
XFILL_35_DFFSR_140 gnd vdd FILL
XFILL_35_DFFSR_151 gnd vdd FILL
XFILL_35_DFFSR_162 gnd vdd FILL
XFILL_35_DFFSR_173 gnd vdd FILL
XFILL_35_DFFSR_184 gnd vdd FILL
XFILL_35_DFFSR_195 gnd vdd FILL
XFILL_1_BUFX4_16 gnd vdd FILL
XFILL_1_BUFX4_27 gnd vdd FILL
XFILL_52_DFFSR_8 gnd vdd FILL
XFILL_7_MUX2X1_130 gnd vdd FILL
XFILL_1_BUFX4_38 gnd vdd FILL
XFILL_7_MUX2X1_141 gnd vdd FILL
XFILL_39_DFFSR_150 gnd vdd FILL
XFILL_1_BUFX4_49 gnd vdd FILL
XFILL_7_MUX2X1_152 gnd vdd FILL
XFILL_39_DFFSR_161 gnd vdd FILL
XFILL_7_MUX2X1_163 gnd vdd FILL
XFILL_39_DFFSR_172 gnd vdd FILL
XFILL_7_MUX2X1_174 gnd vdd FILL
XFILL_7_MUX2X1_185 gnd vdd FILL
XFILL_39_DFFSR_183 gnd vdd FILL
XFILL_39_DFFSR_194 gnd vdd FILL
XFILL_31_NOR3X1_30 gnd vdd FILL
XFILL_13_DFFSR_108 gnd vdd FILL
XFILL_13_DFFSR_119 gnd vdd FILL
XFILL_31_NOR3X1_41 gnd vdd FILL
XFILL_31_NOR3X1_52 gnd vdd FILL
XFILL_58_DFFSR_19 gnd vdd FILL
XNOR2X1_7 NOR2X1_7/A NOR2X1_7/B gnd NOR2X1_9/B vdd NOR2X1
XFILL_81_DFFSR_230 gnd vdd FILL
XFILL_81_DFFSR_241 gnd vdd FILL
XFILL_81_DFFSR_252 gnd vdd FILL
XFILL_81_DFFSR_263 gnd vdd FILL
XFILL_81_DFFSR_274 gnd vdd FILL
XFILL_17_DFFSR_107 gnd vdd FILL
XFILL_17_DFFSR_118 gnd vdd FILL
XFILL_17_DFFSR_129 gnd vdd FILL
XFILL_12_AOI21X1_3 gnd vdd FILL
XFILL_7_INVX1_1 gnd vdd FILL
XFILL_85_DFFSR_240 gnd vdd FILL
XFILL_85_DFFSR_251 gnd vdd FILL
XFILL_85_DFFSR_262 gnd vdd FILL
XFILL_85_DFFSR_273 gnd vdd FILL
XFILL_27_DFFSR_18 gnd vdd FILL
XFILL_66_4 gnd vdd FILL
XFILL_27_DFFSR_29 gnd vdd FILL
XFILL_59_3 gnd vdd FILL
XFILL_1_INVX1_190 gnd vdd FILL
XFILL_8_NAND3X1_120 gnd vdd FILL
XFILL_13_NOR3X1_19 gnd vdd FILL
XFILL_67_DFFSR_17 gnd vdd FILL
XFILL_8_NAND3X1_131 gnd vdd FILL
XFILL_67_DFFSR_28 gnd vdd FILL
XFILL_67_DFFSR_39 gnd vdd FILL
XFILL_63_DFFSR_208 gnd vdd FILL
XFILL_35_4_1 gnd vdd FILL
XFILL_63_DFFSR_219 gnd vdd FILL
XFILL_17_NOR3X1_18 gnd vdd FILL
XFILL_17_NOR3X1_29 gnd vdd FILL
XFILL_67_DFFSR_207 gnd vdd FILL
XFILL_36_DFFSR_16 gnd vdd FILL
XFILL_67_DFFSR_218 gnd vdd FILL
XFILL_67_DFFSR_229 gnd vdd FILL
XFILL_36_DFFSR_27 gnd vdd FILL
XFILL_36_DFFSR_38 gnd vdd FILL
XFILL_36_DFFSR_49 gnd vdd FILL
XAOI21X1_17 BUFX4_80/Y NOR2X1_161/B NOR2X1_158/Y gnd DFFSR_81/D vdd AOI21X1
XAOI21X1_28 BUFX4_65/Y MUX2X1_16/S NOR2X1_183/Y gnd DFFSR_25/D vdd AOI21X1
XFILL_76_DFFSR_15 gnd vdd FILL
XAOI21X1_39 BUFX4_85/Y NOR2X1_202/B NOR2X1_199/Y gnd DFFSR_6/D vdd AOI21X1
XFILL_76_DFFSR_26 gnd vdd FILL
XFILL_76_DFFSR_37 gnd vdd FILL
XFILL_19_MUX2X1_5 gnd vdd FILL
XFILL_76_DFFSR_48 gnd vdd FILL
XFILL_3_NAND2X1_13 gnd vdd FILL
XFILL_3_NAND2X1_24 gnd vdd FILL
XFILL_76_DFFSR_59 gnd vdd FILL
XFILL_3_NAND2X1_35 gnd vdd FILL
XFILL_3_NAND2X1_46 gnd vdd FILL
XFILL_3_NAND2X1_57 gnd vdd FILL
XFILL_3_NAND2X1_68 gnd vdd FILL
XFILL_3_NAND2X1_79 gnd vdd FILL
XFILL_0_AND2X2_3 gnd vdd FILL
XFILL_45_DFFSR_14 gnd vdd FILL
XFILL_45_DFFSR_25 gnd vdd FILL
XFILL_45_DFFSR_36 gnd vdd FILL
XFILL_45_DFFSR_47 gnd vdd FILL
XFILL_45_DFFSR_58 gnd vdd FILL
XFILL_45_DFFSR_69 gnd vdd FILL
XFILL_52_DFFSR_240 gnd vdd FILL
XFILL_85_DFFSR_13 gnd vdd FILL
XFILL_52_DFFSR_251 gnd vdd FILL
XFILL_85_DFFSR_24 gnd vdd FILL
XFILL_52_DFFSR_262 gnd vdd FILL
XFILL_85_DFFSR_35 gnd vdd FILL
XFILL_52_DFFSR_273 gnd vdd FILL
XFILL_12_DFFSR_1 gnd vdd FILL
XFILL_85_DFFSR_46 gnd vdd FILL
XFILL_29_CLKBUF1_12 gnd vdd FILL
XFILL_14_DFFSR_13 gnd vdd FILL
XFILL_85_DFFSR_57 gnd vdd FILL
XFILL_29_CLKBUF1_23 gnd vdd FILL
XFILL_85_DFFSR_68 gnd vdd FILL
XFILL_14_DFFSR_24 gnd vdd FILL
XFILL_14_DFFSR_35 gnd vdd FILL
XFILL_29_CLKBUF1_34 gnd vdd FILL
XFILL_85_DFFSR_79 gnd vdd FILL
XFILL_14_DFFSR_46 gnd vdd FILL
XFILL_14_DFFSR_57 gnd vdd FILL
XFILL_26_4_1 gnd vdd FILL
XFILL_56_DFFSR_250 gnd vdd FILL
XFILL_14_DFFSR_68 gnd vdd FILL
XFILL_3_AOI22X1_11 gnd vdd FILL
XFILL_1_4_1 gnd vdd FILL
XFILL_56_DFFSR_261 gnd vdd FILL
XFILL_56_DFFSR_272 gnd vdd FILL
XFILL_14_DFFSR_79 gnd vdd FILL
XFILL_11_CLKBUF1_2 gnd vdd FILL
XFILL_30_DFFSR_208 gnd vdd FILL
XFILL_54_DFFSR_12 gnd vdd FILL
XFILL_7_AOI21X1_13 gnd vdd FILL
XFILL_30_DFFSR_219 gnd vdd FILL
XOAI22X1_14 INVX1_41/Y INVX1_121/A INVX1_43/Y INVX1_120/A gnd NOR3X1_20/C vdd OAI22X1
XFILL_54_DFFSR_23 gnd vdd FILL
XFILL_7_AOI21X1_24 gnd vdd FILL
XFILL_54_DFFSR_34 gnd vdd FILL
XOAI22X1_25 INVX1_186/Y OAI22X1_50/B INVX1_181/Y OAI22X1_50/D gnd NOR2X1_83/B vdd
+ OAI22X1
XFILL_25_NOR3X1_9 gnd vdd FILL
XFILL_7_AOI21X1_35 gnd vdd FILL
XFILL_54_DFFSR_45 gnd vdd FILL
XFILL_54_DFFSR_56 gnd vdd FILL
XFILL_83_DFFSR_150 gnd vdd FILL
XOAI22X1_36 INVX1_29/Y OAI22X1_36/B MUX2X1_3/B OAI22X1_36/D gnd NOR2X1_97/B vdd OAI22X1
XFILL_83_DFFSR_161 gnd vdd FILL
XFILL_7_AOI21X1_46 gnd vdd FILL
XOAI22X1_47 INVX1_132/A INVX1_130/Y INVX1_131/Y INVX1_133/A gnd AOI22X1_3/A vdd OAI22X1
XFILL_54_DFFSR_67 gnd vdd FILL
XFILL_17_OAI22X1_15 gnd vdd FILL
XFILL_7_AOI21X1_57 gnd vdd FILL
XFILL_54_DFFSR_78 gnd vdd FILL
XFILL_7_AOI21X1_68 gnd vdd FILL
XFILL_15_CLKBUF1_1 gnd vdd FILL
XFILL_83_DFFSR_172 gnd vdd FILL
XFILL_54_DFFSR_89 gnd vdd FILL
XFILL_83_DFFSR_183 gnd vdd FILL
XFILL_17_OAI22X1_26 gnd vdd FILL
XFILL_7_AOI21X1_79 gnd vdd FILL
XFILL_83_DFFSR_194 gnd vdd FILL
XFILL_17_OAI22X1_37 gnd vdd FILL
XFILL_34_DFFSR_207 gnd vdd FILL
XFILL_3_DFFSR_220 gnd vdd FILL
XFILL_17_OAI22X1_48 gnd vdd FILL
XFILL_34_DFFSR_218 gnd vdd FILL
XFILL_3_DFFSR_231 gnd vdd FILL
XFILL_34_DFFSR_229 gnd vdd FILL
XFILL_3_DFFSR_242 gnd vdd FILL
XFILL_34_DFFSR_5 gnd vdd FILL
XFILL_23_DFFSR_11 gnd vdd FILL
XFILL_3_DFFSR_253 gnd vdd FILL
XFILL_87_DFFSR_160 gnd vdd FILL
XFILL_3_DFFSR_264 gnd vdd FILL
XFILL_3_DFFSR_275 gnd vdd FILL
XFILL_1_CLKBUF1_16 gnd vdd FILL
XFILL_23_DFFSR_22 gnd vdd FILL
XFILL_87_DFFSR_171 gnd vdd FILL
XFILL_23_DFFSR_33 gnd vdd FILL
XFILL_1_CLKBUF1_27 gnd vdd FILL
XFILL_87_DFFSR_182 gnd vdd FILL
XFILL_23_DFFSR_44 gnd vdd FILL
XFILL_1_CLKBUF1_38 gnd vdd FILL
XFILL_61_DFFSR_107 gnd vdd FILL
XFILL_23_DFFSR_55 gnd vdd FILL
XFILL_87_DFFSR_193 gnd vdd FILL
XFILL_38_DFFSR_206 gnd vdd FILL
XFILL_23_DFFSR_66 gnd vdd FILL
XFILL_38_DFFSR_217 gnd vdd FILL
XFILL_7_DFFSR_230 gnd vdd FILL
XFILL_61_DFFSR_118 gnd vdd FILL
XFILL_23_DFFSR_77 gnd vdd FILL
XFILL_38_DFFSR_228 gnd vdd FILL
XFILL_61_DFFSR_129 gnd vdd FILL
XFILL_7_DFFSR_241 gnd vdd FILL
XFILL_23_DFFSR_88 gnd vdd FILL
XFILL_23_DFFSR_99 gnd vdd FILL
XFILL_38_DFFSR_239 gnd vdd FILL
XFILL_7_DFFSR_252 gnd vdd FILL
XFILL_63_DFFSR_10 gnd vdd FILL
XFILL_63_DFFSR_21 gnd vdd FILL
XFILL_7_DFFSR_263 gnd vdd FILL
XFILL_7_DFFSR_274 gnd vdd FILL
XFILL_63_DFFSR_32 gnd vdd FILL
XFILL_63_DFFSR_43 gnd vdd FILL
XFILL_4_MUX2X1_19 gnd vdd FILL
XFILL_65_DFFSR_106 gnd vdd FILL
XFILL_63_DFFSR_54 gnd vdd FILL
XFILL_63_DFFSR_65 gnd vdd FILL
XFILL_63_DFFSR_76 gnd vdd FILL
XFILL_10_OAI21X1_17 gnd vdd FILL
XFILL_65_DFFSR_117 gnd vdd FILL
XFILL_10_OAI21X1_28 gnd vdd FILL
XFILL_9_5_1 gnd vdd FILL
XFILL_65_DFFSR_128 gnd vdd FILL
XFILL_63_DFFSR_87 gnd vdd FILL
XFILL_10_OAI21X1_39 gnd vdd FILL
XFILL_65_DFFSR_139 gnd vdd FILL
XFILL_63_DFFSR_98 gnd vdd FILL
XFILL_8_0_0 gnd vdd FILL
XFILL_6_DFFSR_12 gnd vdd FILL
XFILL_8_MUX2X1_18 gnd vdd FILL
XFILL_6_DFFSR_23 gnd vdd FILL
XFILL_69_DFFSR_105 gnd vdd FILL
XFILL_8_MUX2X1_29 gnd vdd FILL
XFILL_6_DFFSR_34 gnd vdd FILL
XFILL_32_DFFSR_20 gnd vdd FILL
XFILL_69_DFFSR_116 gnd vdd FILL
XFILL_6_DFFSR_45 gnd vdd FILL
XFILL_56_DFFSR_9 gnd vdd FILL
XFILL_6_DFFSR_56 gnd vdd FILL
XFILL_32_DFFSR_31 gnd vdd FILL
XFILL_6_DFFSR_67 gnd vdd FILL
XFILL_69_DFFSR_127 gnd vdd FILL
XFILL_69_DFFSR_138 gnd vdd FILL
XFILL_32_DFFSR_42 gnd vdd FILL
XFILL_0_AOI22X1_3 gnd vdd FILL
XFILL_69_DFFSR_149 gnd vdd FILL
XFILL_6_DFFSR_78 gnd vdd FILL
XFILL_12_OAI21X1_6 gnd vdd FILL
XFILL_32_DFFSR_53 gnd vdd FILL
XFILL_7_OAI22X1_10 gnd vdd FILL
XFILL_6_DFFSR_89 gnd vdd FILL
XFILL_32_DFFSR_64 gnd vdd FILL
XFILL_7_OAI22X1_21 gnd vdd FILL
XFILL_32_DFFSR_75 gnd vdd FILL
XFILL_7_OAI22X1_32 gnd vdd FILL
XFILL_32_DFFSR_86 gnd vdd FILL
XFILL_7_OAI22X1_43 gnd vdd FILL
XFILL_0_INVX1_202 gnd vdd FILL
XFILL_32_DFFSR_97 gnd vdd FILL
XFILL_0_INVX1_213 gnd vdd FILL
XFILL_72_DFFSR_30 gnd vdd FILL
XFILL_0_INVX1_224 gnd vdd FILL
XFILL_72_DFFSR_41 gnd vdd FILL
XFILL_17_4_1 gnd vdd FILL
XFILL_4_AOI22X1_2 gnd vdd FILL
XFILL_72_DFFSR_52 gnd vdd FILL
XFILL_72_DFFSR_63 gnd vdd FILL
XFILL_72_DFFSR_74 gnd vdd FILL
XFILL_23_DFFSR_250 gnd vdd FILL
XFILL_72_DFFSR_85 gnd vdd FILL
XFILL_23_DFFSR_261 gnd vdd FILL
XFILL_23_DFFSR_272 gnd vdd FILL
XFILL_72_DFFSR_96 gnd vdd FILL
XFILL_60_7_2 gnd vdd FILL
XFILL_4_INVX1_201 gnd vdd FILL
XFILL_4_INVX1_212 gnd vdd FILL
XFILL_20_MUX2X1_17 gnd vdd FILL
XFILL_4_INVX1_223 gnd vdd FILL
XFILL_20_MUX2X1_28 gnd vdd FILL
XFILL_4_NOR2X1_201 gnd vdd FILL
XFILL_20_MUX2X1_39 gnd vdd FILL
XFILL_8_AOI22X1_1 gnd vdd FILL
XFILL_50_DFFSR_150 gnd vdd FILL
XFILL_50_DFFSR_161 gnd vdd FILL
XFILL_41_DFFSR_40 gnd vdd FILL
XFILL_27_DFFSR_260 gnd vdd FILL
XFILL_12_NOR3X1_4 gnd vdd FILL
XFILL_27_DFFSR_271 gnd vdd FILL
XFILL_41_DFFSR_51 gnd vdd FILL
XFILL_50_DFFSR_172 gnd vdd FILL
XFILL_0_OAI21X1_12 gnd vdd FILL
XFILL_50_DFFSR_183 gnd vdd FILL
XFILL_50_DFFSR_194 gnd vdd FILL
XFILL_41_DFFSR_62 gnd vdd FILL
XFILL_0_OAI21X1_23 gnd vdd FILL
XFILL_41_DFFSR_73 gnd vdd FILL
XFILL_0_OAI21X1_34 gnd vdd FILL
XFILL_41_DFFSR_84 gnd vdd FILL
XFILL_0_OAI21X1_45 gnd vdd FILL
XFILL_18_CLKBUF1_30 gnd vdd FILL
XFILL_41_DFFSR_95 gnd vdd FILL
XFILL_18_CLKBUF1_41 gnd vdd FILL
XFILL_54_DFFSR_160 gnd vdd FILL
XFILL_54_DFFSR_171 gnd vdd FILL
XFILL_81_DFFSR_50 gnd vdd FILL
XFILL_81_DFFSR_61 gnd vdd FILL
XFILL_54_DFFSR_182 gnd vdd FILL
XFILL_54_DFFSR_193 gnd vdd FILL
XFILL_13_AOI21X1_60 gnd vdd FILL
XFILL_13_AOI21X1_71 gnd vdd FILL
XFILL_81_DFFSR_72 gnd vdd FILL
XFILL_81_DFFSR_83 gnd vdd FILL
XFILL_81_DFFSR_94 gnd vdd FILL
XFILL_10_DFFSR_50 gnd vdd FILL
XFILL_10_DFFSR_61 gnd vdd FILL
XFILL_10_DFFSR_72 gnd vdd FILL
XFILL_10_DFFSR_83 gnd vdd FILL
XFILL_58_DFFSR_170 gnd vdd FILL
XFILL_10_DFFSR_94 gnd vdd FILL
XFILL_58_DFFSR_181 gnd vdd FILL
XFILL_32_DFFSR_106 gnd vdd FILL
XFILL_58_DFFSR_192 gnd vdd FILL
XFILL_21_NOR3X1_2 gnd vdd FILL
XFILL_1_DFFSR_130 gnd vdd FILL
XFILL_32_DFFSR_117 gnd vdd FILL
XFILL_32_DFFSR_128 gnd vdd FILL
XFILL_1_DFFSR_141 gnd vdd FILL
XFILL_1_DFFSR_152 gnd vdd FILL
XFILL_50_DFFSR_60 gnd vdd FILL
XFILL_32_DFFSR_139 gnd vdd FILL
XFILL_1_DFFSR_163 gnd vdd FILL
XFILL_50_DFFSR_71 gnd vdd FILL
XFILL_21_13 gnd vdd FILL
XFILL_50_DFFSR_82 gnd vdd FILL
XFILL_1_DFFSR_174 gnd vdd FILL
XFILL_50_DFFSR_93 gnd vdd FILL
XFILL_1_DFFSR_185 gnd vdd FILL
XFILL_1_DFFSR_196 gnd vdd FILL
XFILL_36_DFFSR_105 gnd vdd FILL
XFILL_36_DFFSR_116 gnd vdd FILL
XFILL_5_DFFSR_140 gnd vdd FILL
XFILL_36_DFFSR_127 gnd vdd FILL
XFILL_36_DFFSR_138 gnd vdd FILL
XFILL_5_DFFSR_151 gnd vdd FILL
XFILL_5_DFFSR_162 gnd vdd FILL
XFILL_36_DFFSR_149 gnd vdd FILL
XFILL_5_DFFSR_173 gnd vdd FILL
XFILL_5_DFFSR_184 gnd vdd FILL
XFILL_9_NAND3X1_110 gnd vdd FILL
XFILL_9_NAND3X1_121 gnd vdd FILL
XFILL_5_DFFSR_195 gnd vdd FILL
XFILL_9_NAND3X1_132 gnd vdd FILL
XFILL_16_MUX2X1_110 gnd vdd FILL
XFILL_16_MUX2X1_121 gnd vdd FILL
XFILL_4_NOR3X1_3 gnd vdd FILL
XFILL_9_DFFSR_150 gnd vdd FILL
XFILL_9_DFFSR_161 gnd vdd FILL
XFILL_51_7_2 gnd vdd FILL
XFILL_9_DFFSR_172 gnd vdd FILL
XFILL_13_MUX2X1_70 gnd vdd FILL
XFILL_16_MUX2X1_132 gnd vdd FILL
XFILL_16_MUX2X1_143 gnd vdd FILL
XFILL_13_MUX2X1_81 gnd vdd FILL
XFILL_50_2_1 gnd vdd FILL
XFILL_16_MUX2X1_154 gnd vdd FILL
XFILL_9_DFFSR_183 gnd vdd FILL
XFILL_16_MUX2X1_165 gnd vdd FILL
XFILL_13_MUX2X1_92 gnd vdd FILL
XFILL_9_DFFSR_194 gnd vdd FILL
XFILL_1_NOR3X1_30 gnd vdd FILL
XFILL_1_NOR3X1_41 gnd vdd FILL
XFILL_16_MUX2X1_176 gnd vdd FILL
XFILL_16_MUX2X1_187 gnd vdd FILL
XFILL_1_NOR3X1_52 gnd vdd FILL
XFILL_82_DFFSR_206 gnd vdd FILL
XFILL_82_DFFSR_217 gnd vdd FILL
XFILL_82_DFFSR_228 gnd vdd FILL
XFILL_17_MUX2X1_80 gnd vdd FILL
XFILL_3_DFFSR_4 gnd vdd FILL
XFILL_82_DFFSR_239 gnd vdd FILL
XFILL_17_MUX2X1_91 gnd vdd FILL
XFILL_16_DFFSR_2 gnd vdd FILL
XFILL_5_NOR3X1_40 gnd vdd FILL
XFILL_73_DFFSR_3 gnd vdd FILL
XFILL_5_NOR3X1_51 gnd vdd FILL
XFILL_2_DFFSR_60 gnd vdd FILL
XFILL_2_DFFSR_71 gnd vdd FILL
XFILL_2_DFFSR_82 gnd vdd FILL
XFILL_86_DFFSR_205 gnd vdd FILL
XFILL_86_DFFSR_216 gnd vdd FILL
XFILL_2_DFFSR_93 gnd vdd FILL
XFILL_86_DFFSR_227 gnd vdd FILL
XFILL_86_DFFSR_238 gnd vdd FILL
XFILL_21_DFFSR_160 gnd vdd FILL
XFILL_86_DFFSR_249 gnd vdd FILL
XFILL_2_INVX1_100 gnd vdd FILL
XFILL_21_DFFSR_171 gnd vdd FILL
XFILL_2_INVX1_111 gnd vdd FILL
XFILL_21_DFFSR_182 gnd vdd FILL
XFILL_9_NOR3X1_50 gnd vdd FILL
XFILL_21_DFFSR_193 gnd vdd FILL
XFILL_11_BUFX2_8 gnd vdd FILL
XFILL_2_INVX1_122 gnd vdd FILL
XFILL_2_INVX1_133 gnd vdd FILL
XFILL_2_INVX1_144 gnd vdd FILL
XFILL_2_INVX1_155 gnd vdd FILL
XFILL_2_INVX1_166 gnd vdd FILL
XFILL_25_DFFSR_170 gnd vdd FILL
XFILL_2_INVX1_177 gnd vdd FILL
XFILL_2_INVX1_188 gnd vdd FILL
XFILL_2_INVX1_199 gnd vdd FILL
XFILL_6_INVX1_110 gnd vdd FILL
XFILL_25_DFFSR_181 gnd vdd FILL
XFILL_6_INVX1_121 gnd vdd FILL
XFILL_25_DFFSR_192 gnd vdd FILL
XFILL_6_INVX1_132 gnd vdd FILL
XFILL_58_3_1 gnd vdd FILL
XFILL_6_INVX1_143 gnd vdd FILL
XFILL_6_INVX1_154 gnd vdd FILL
XFILL_6_INVX1_165 gnd vdd FILL
XFILL_38_DFFSR_6 gnd vdd FILL
XFILL_6_MUX2X1_160 gnd vdd FILL
XFILL_6_MUX2X1_171 gnd vdd FILL
XFILL_6_INVX1_176 gnd vdd FILL
XFILL_29_DFFSR_180 gnd vdd FILL
XFILL_6_INVX1_187 gnd vdd FILL
XFILL_6_MUX2X1_182 gnd vdd FILL
XFILL_6_INVX1_198 gnd vdd FILL
XFILL_6_MUX2X1_193 gnd vdd FILL
XFILL_29_DFFSR_191 gnd vdd FILL
XFILL_0_OAI22X1_6 gnd vdd FILL
XFILL_71_DFFSR_260 gnd vdd FILL
XFILL_71_DFFSR_271 gnd vdd FILL
XFILL_42_7_2 gnd vdd FILL
XFILL_41_2_1 gnd vdd FILL
XFILL_4_OAI22X1_5 gnd vdd FILL
XFILL_10_BUFX4_2 gnd vdd FILL
XFILL_75_DFFSR_270 gnd vdd FILL
XFILL_8_OAI22X1_4 gnd vdd FILL
XFILL_53_DFFSR_205 gnd vdd FILL
XFILL_53_DFFSR_216 gnd vdd FILL
XFILL_53_DFFSR_227 gnd vdd FILL
XFILL_9_NAND3X1_30 gnd vdd FILL
XFILL_53_DFFSR_238 gnd vdd FILL
XFILL_9_NAND3X1_41 gnd vdd FILL
XFILL_53_DFFSR_249 gnd vdd FILL
XFILL_9_NAND3X1_52 gnd vdd FILL
XFILL_9_NAND3X1_63 gnd vdd FILL
XFILL_15_BUFX4_10 gnd vdd FILL
XFILL_9_NAND3X1_74 gnd vdd FILL
XFILL_15_BUFX4_21 gnd vdd FILL
XFILL_80_DFFSR_105 gnd vdd FILL
XFILL_9_NAND3X1_85 gnd vdd FILL
XFILL_15_BUFX4_32 gnd vdd FILL
XFILL_9_NAND3X1_96 gnd vdd FILL
XFILL_57_DFFSR_204 gnd vdd FILL
XFILL_57_DFFSR_215 gnd vdd FILL
XFILL_15_BUFX4_43 gnd vdd FILL
XFILL_80_DFFSR_116 gnd vdd FILL
XFILL_15_BUFX4_54 gnd vdd FILL
XFILL_80_DFFSR_127 gnd vdd FILL
XFILL_57_DFFSR_226 gnd vdd FILL
XFILL_80_DFFSR_138 gnd vdd FILL
XFILL_57_DFFSR_237 gnd vdd FILL
XFILL_15_BUFX4_65 gnd vdd FILL
XFILL_80_DFFSR_149 gnd vdd FILL
XFILL_15_BUFX4_76 gnd vdd FILL
XFILL_57_DFFSR_248 gnd vdd FILL
XFILL_15_BUFX4_87 gnd vdd FILL
XFILL_49_3_1 gnd vdd FILL
XFILL_57_DFFSR_259 gnd vdd FILL
XFILL_15_BUFX4_98 gnd vdd FILL
XFILL_84_DFFSR_104 gnd vdd FILL
XFILL_0_DFFSR_208 gnd vdd FILL
XFILL_0_DFFSR_219 gnd vdd FILL
XFILL_84_DFFSR_115 gnd vdd FILL
XFILL_84_DFFSR_126 gnd vdd FILL
XFILL_84_DFFSR_137 gnd vdd FILL
XFILL_84_DFFSR_148 gnd vdd FILL
XFILL_2_NAND2X1_10 gnd vdd FILL
XFILL_84_DFFSR_159 gnd vdd FILL
XFILL_2_NAND2X1_21 gnd vdd FILL
XFILL_2_NAND2X1_32 gnd vdd FILL
XFILL_4_DFFSR_207 gnd vdd FILL
XFILL_2_NAND2X1_43 gnd vdd FILL
XFILL_1_NAND3X1_7 gnd vdd FILL
XFILL_4_DFFSR_218 gnd vdd FILL
XFILL_2_NAND2X1_54 gnd vdd FILL
XFILL_2_NAND2X1_65 gnd vdd FILL
XFILL_4_DFFSR_229 gnd vdd FILL
XFILL_0_INVX8_2 gnd vdd FILL
XFILL_2_NAND2X1_76 gnd vdd FILL
XFILL_2_NAND2X1_87 gnd vdd FILL
XFILL_33_7_2 gnd vdd FILL
XFILL_12_BUFX4_105 gnd vdd FILL
XFILL_32_2_1 gnd vdd FILL
XFILL_8_DFFSR_206 gnd vdd FILL
XFILL_10_CLKBUF1_18 gnd vdd FILL
XFILL_5_NAND3X1_6 gnd vdd FILL
XFILL_8_DFFSR_217 gnd vdd FILL
XFILL_10_CLKBUF1_29 gnd vdd FILL
XFILL_8_DFFSR_228 gnd vdd FILL
XFILL_8_DFFSR_239 gnd vdd FILL
XFILL_73_DFFSR_19 gnd vdd FILL
XFILL_42_DFFSR_270 gnd vdd FILL
XFILL_9_NAND3X1_5 gnd vdd FILL
XFILL_16_MUX2X1_9 gnd vdd FILL
XFILL_28_CLKBUF1_20 gnd vdd FILL
XFILL_16_13 gnd vdd FILL
XFILL_28_CLKBUF1_31 gnd vdd FILL
XFILL_28_CLKBUF1_42 gnd vdd FILL
XFILL_7_BUFX4_20 gnd vdd FILL
XFILL_7_BUFX4_31 gnd vdd FILL
XFILL_7_BUFX4_42 gnd vdd FILL
XFILL_7_BUFX4_53 gnd vdd FILL
XFILL_7_BUFX4_64 gnd vdd FILL
XFILL_42_DFFSR_18 gnd vdd FILL
XFILL_20_DFFSR_205 gnd vdd FILL
XFILL_42_DFFSR_29 gnd vdd FILL
XFILL_7_BUFX4_75 gnd vdd FILL
XFILL_19_MUX2X1_109 gnd vdd FILL
XFILL_6_AOI21X1_10 gnd vdd FILL
XFILL_20_DFFSR_216 gnd vdd FILL
XFILL_7_BUFX4_86 gnd vdd FILL
XFILL_10_NOR2X1_18 gnd vdd FILL
XFILL_7_BUFX4_97 gnd vdd FILL
XFILL_6_AOI21X1_21 gnd vdd FILL
XFILL_20_DFFSR_227 gnd vdd FILL
XFILL_10_NOR2X1_29 gnd vdd FILL
XFILL_6_AOI21X1_32 gnd vdd FILL
XFILL_20_DFFSR_238 gnd vdd FILL
XFILL_6_AOI21X1_43 gnd vdd FILL
XFILL_20_DFFSR_249 gnd vdd FILL
XFILL_6_AOI21X1_54 gnd vdd FILL
XFILL_16_OAI22X1_12 gnd vdd FILL
XFILL_16_OAI22X1_23 gnd vdd FILL
XFILL_6_AOI21X1_65 gnd vdd FILL
XFILL_73_DFFSR_180 gnd vdd FILL
XFILL_6_AOI21X1_76 gnd vdd FILL
XFILL_82_DFFSR_17 gnd vdd FILL
XFILL_16_OAI22X1_34 gnd vdd FILL
XFILL_73_DFFSR_191 gnd vdd FILL
XFILL_82_DFFSR_28 gnd vdd FILL
XFILL_24_DFFSR_204 gnd vdd FILL
XFILL_16_OAI22X1_45 gnd vdd FILL
XFILL_24_DFFSR_215 gnd vdd FILL
XFILL_82_DFFSR_39 gnd vdd FILL
XFILL_24_DFFSR_226 gnd vdd FILL
XFILL_9_NOR2X1_120 gnd vdd FILL
XFILL_9_NOR2X1_131 gnd vdd FILL
XFILL_7_DFFSR_5 gnd vdd FILL
XFILL_24_DFFSR_237 gnd vdd FILL
XFILL_11_DFFSR_17 gnd vdd FILL
XFILL_24_DFFSR_248 gnd vdd FILL
XFILL_11_DFFSR_28 gnd vdd FILL
XFILL_9_NOR2X1_142 gnd vdd FILL
XFILL_9_NOR2X1_153 gnd vdd FILL
XFILL_11_DFFSR_39 gnd vdd FILL
XFILL_0_CLKBUF1_13 gnd vdd FILL
XFILL_24_DFFSR_259 gnd vdd FILL
XFILL_0_CLKBUF1_24 gnd vdd FILL
XFILL_9_NOR2X1_164 gnd vdd FILL
XFILL_77_DFFSR_4 gnd vdd FILL
XFILL_9_NOR2X1_175 gnd vdd FILL
XFILL_0_CLKBUF1_35 gnd vdd FILL
XFILL_51_DFFSR_104 gnd vdd FILL
XFILL_77_DFFSR_190 gnd vdd FILL
XFILL_28_DFFSR_203 gnd vdd FILL
XFILL_9_NOR2X1_186 gnd vdd FILL
XFILL_9_NOR2X1_197 gnd vdd FILL
XFILL_51_DFFSR_115 gnd vdd FILL
XFILL_28_DFFSR_214 gnd vdd FILL
XFILL_51_DFFSR_126 gnd vdd FILL
XFILL_28_DFFSR_225 gnd vdd FILL
XFILL_51_DFFSR_137 gnd vdd FILL
XFILL_28_DFFSR_236 gnd vdd FILL
XFILL_51_DFFSR_148 gnd vdd FILL
XFILL_51_DFFSR_16 gnd vdd FILL
XFILL_28_DFFSR_247 gnd vdd FILL
XFILL_51_DFFSR_27 gnd vdd FILL
XFILL_51_DFFSR_159 gnd vdd FILL
XFILL_51_DFFSR_38 gnd vdd FILL
XFILL_28_DFFSR_258 gnd vdd FILL
XFILL_28_DFFSR_269 gnd vdd FILL
XFILL_51_DFFSR_49 gnd vdd FILL
XFILL_55_DFFSR_103 gnd vdd FILL
XFILL_24_7_2 gnd vdd FILL
XFILL_55_DFFSR_114 gnd vdd FILL
XFILL_23_2_1 gnd vdd FILL
XFILL_55_DFFSR_125 gnd vdd FILL
XFILL_55_DFFSR_136 gnd vdd FILL
XFILL_55_DFFSR_147 gnd vdd FILL
XFILL_55_DFFSR_158 gnd vdd FILL
XFILL_8_MUX2X1_8 gnd vdd FILL
XFILL_55_DFFSR_169 gnd vdd FILL
XFILL_20_DFFSR_15 gnd vdd FILL
XFILL_59_DFFSR_102 gnd vdd FILL
XFILL_9_MUX2X1_104 gnd vdd FILL
XFILL_9_MUX2X1_115 gnd vdd FILL
XFILL_20_DFFSR_26 gnd vdd FILL
XFILL_59_DFFSR_113 gnd vdd FILL
XFILL_59_DFFSR_124 gnd vdd FILL
XFILL_20_DFFSR_37 gnd vdd FILL
XFILL_9_MUX2X1_126 gnd vdd FILL
XFILL_20_DFFSR_48 gnd vdd FILL
XFILL_9_MUX2X1_137 gnd vdd FILL
XFILL_11_BUFX4_80 gnd vdd FILL
XFILL_59_DFFSR_135 gnd vdd FILL
XFILL_20_DFFSR_59 gnd vdd FILL
XFILL_59_DFFSR_146 gnd vdd FILL
XFILL_11_BUFX4_91 gnd vdd FILL
XFILL_9_MUX2X1_148 gnd vdd FILL
XFILL_59_DFFSR_157 gnd vdd FILL
XFILL_9_MUX2X1_159 gnd vdd FILL
XFILL_59_DFFSR_168 gnd vdd FILL
XFILL_59_DFFSR_179 gnd vdd FILL
XFILL_6_OAI22X1_40 gnd vdd FILL
XFILL_2_DFFSR_106 gnd vdd FILL
XFILL_60_DFFSR_14 gnd vdd FILL
XFILL_6_OAI22X1_51 gnd vdd FILL
XFILL_60_DFFSR_25 gnd vdd FILL
XFILL_2_DFFSR_117 gnd vdd FILL
XFILL_60_DFFSR_36 gnd vdd FILL
XFILL_2_DFFSR_128 gnd vdd FILL
XFILL_2_DFFSR_139 gnd vdd FILL
XDFFSR_50 INVX1_7/A DFFSR_76/CLK DFFSR_53/R vdd DFFSR_50/D gnd vdd DFFSR
XFILL_60_DFFSR_47 gnd vdd FILL
XFILL_60_DFFSR_58 gnd vdd FILL
XDFFSR_61 DFFSR_61/Q DFFSR_97/CLK DFFSR_69/R vdd DFFSR_61/D gnd vdd DFFSR
XFILL_60_DFFSR_69 gnd vdd FILL
XDFFSR_72 DFFSR_72/Q DFFSR_72/CLK DFFSR_96/R vdd DFFSR_72/D gnd vdd DFFSR
XDFFSR_83 DFFSR_83/Q DFFSR_84/CLK DFFSR_84/R vdd DFFSR_83/D gnd vdd DFFSR
XDFFSR_94 DFFSR_94/Q DFFSR_94/CLK DFFSR_99/R vdd DFFSR_94/D gnd vdd DFFSR
XFILL_6_DFFSR_105 gnd vdd FILL
XFILL_6_DFFSR_116 gnd vdd FILL
XFILL_10_MUX2X1_14 gnd vdd FILL
XFILL_3_DFFSR_16 gnd vdd FILL
XFILL_10_MUX2X1_25 gnd vdd FILL
XFILL_6_DFFSR_127 gnd vdd FILL
XFILL_6_DFFSR_138 gnd vdd FILL
XFILL_3_DFFSR_27 gnd vdd FILL
XFILL_10_MUX2X1_36 gnd vdd FILL
XFILL_6_DFFSR_149 gnd vdd FILL
XFILL_3_DFFSR_38 gnd vdd FILL
XFILL_10_MUX2X1_47 gnd vdd FILL
XFILL_1_BUFX4_5 gnd vdd FILL
XFILL_1_AOI21X1_1 gnd vdd FILL
XFILL_10_MUX2X1_58 gnd vdd FILL
XFILL_3_DFFSR_49 gnd vdd FILL
XFILL_14_BUFX4_3 gnd vdd FILL
XFILL_10_MUX2X1_69 gnd vdd FILL
XFILL_40_DFFSR_180 gnd vdd FILL
XFILL_14_MUX2X1_13 gnd vdd FILL
XFILL_6_3_1 gnd vdd FILL
XFILL_5_INVX1_70 gnd vdd FILL
XFILL_40_DFFSR_191 gnd vdd FILL
XFILL_14_MUX2X1_24 gnd vdd FILL
XFILL_5_INVX1_81 gnd vdd FILL
XFILL_14_MUX2X1_35 gnd vdd FILL
XFILL_5_INVX1_92 gnd vdd FILL
XFILL_14_MUX2X1_46 gnd vdd FILL
XFILL_14_MUX2X1_57 gnd vdd FILL
XFILL_14_MUX2X1_68 gnd vdd FILL
XFILL_14_MUX2X1_79 gnd vdd FILL
XFILL_12_MUX2X1_2 gnd vdd FILL
XFILL_2_NOR3X1_17 gnd vdd FILL
XFILL_2_NOR3X1_28 gnd vdd FILL
XFILL_2_NOR3X1_39 gnd vdd FILL
XFILL_18_MUX2X1_12 gnd vdd FILL
XFILL_18_MUX2X1_23 gnd vdd FILL
XFILL_44_DFFSR_190 gnd vdd FILL
XFILL_18_MUX2X1_34 gnd vdd FILL
XFILL_18_MUX2X1_45 gnd vdd FILL
XFILL_18_MUX2X1_56 gnd vdd FILL
XFILL_0_INVX1_9 gnd vdd FILL
XFILL_18_MUX2X1_67 gnd vdd FILL
XFILL_18_MUX2X1_78 gnd vdd FILL
XFILL_15_7_2 gnd vdd FILL
XFILL_6_NOR3X1_16 gnd vdd FILL
XFILL_6_NOR3X1_27 gnd vdd FILL
XFILL_14_2_1 gnd vdd FILL
XFILL_18_MUX2X1_89 gnd vdd FILL
XFILL_6_NOR3X1_38 gnd vdd FILL
XFILL_6_NOR3X1_49 gnd vdd FILL
XFILL_22_DFFSR_103 gnd vdd FILL
XFILL_3_BUFX4_90 gnd vdd FILL
XFILL_22_DFFSR_114 gnd vdd FILL
XFILL_22_DFFSR_125 gnd vdd FILL
XFILL_22_DFFSR_136 gnd vdd FILL
XFILL_22_DFFSR_147 gnd vdd FILL
XFILL_22_DFFSR_158 gnd vdd FILL
XFILL_22_DFFSR_169 gnd vdd FILL
XFILL_3_INVX1_109 gnd vdd FILL
XFILL_26_DFFSR_102 gnd vdd FILL
XFILL_26_DFFSR_113 gnd vdd FILL
XFILL_26_DFFSR_124 gnd vdd FILL
XFILL_1_NAND3X1_18 gnd vdd FILL
XFILL_26_DFFSR_135 gnd vdd FILL
XFILL_1_NAND3X1_29 gnd vdd FILL
XFILL_26_DFFSR_146 gnd vdd FILL
XFILL_26_DFFSR_157 gnd vdd FILL
XINVX1_100 INVX1_100/A gnd MUX2X1_87/A vdd INVX1
XFILL_26_DFFSR_168 gnd vdd FILL
XINVX1_111 DFFSR_79/Q gnd MUX2X1_98/A vdd INVX1
XFILL_5_NOR2X1_3 gnd vdd FILL
XFILL_26_DFFSR_179 gnd vdd FILL
XFILL_7_INVX1_108 gnd vdd FILL
XINVX1_122 NOR2X1_80/B gnd INVX1_122/Y vdd INVX1
XINVX1_133 INVX1_133/A gnd INVX1_133/Y vdd INVX1
XFILL_7_INVX1_119 gnd vdd FILL
XINVX1_144 INVX1_144/A gnd MUX2X1_1/B vdd INVX1
XINVX1_155 INVX1_155/A gnd OAI21X1_3/A vdd INVX1
XINVX1_166 INVX1_166/A gnd NOR2X1_10/B vdd INVX1
XFILL_4_INVX8_3 gnd vdd FILL
XINVX1_177 INVX1_177/A gnd INVX1_177/Y vdd INVX1
XINVX1_188 INVX1_188/A gnd OAI21X1_7/A vdd INVX1
XFILL_17_INVX8_1 gnd vdd FILL
XFILL_15_MUX2X1_140 gnd vdd FILL
XFILL_29_DFFSR_70 gnd vdd FILL
XINVX1_199 DFFSR_92/Q gnd INVX1_199/Y vdd INVX1
XFILL_29_DFFSR_81 gnd vdd FILL
XFILL_15_MUX2X1_151 gnd vdd FILL
XFILL_22_NOR3X1_14 gnd vdd FILL
XFILL_15_MUX2X1_162 gnd vdd FILL
XFILL_29_DFFSR_92 gnd vdd FILL
XFILL_15_MUX2X1_173 gnd vdd FILL
XFILL_22_NOR3X1_25 gnd vdd FILL
XFILL_22_NOR3X1_36 gnd vdd FILL
XFILL_22_NOR3X1_47 gnd vdd FILL
XFILL_15_MUX2X1_184 gnd vdd FILL
XFILL_72_DFFSR_203 gnd vdd FILL
XFILL_4_MUX2X1_1 gnd vdd FILL
XFILL_72_DFFSR_214 gnd vdd FILL
XFILL_72_DFFSR_225 gnd vdd FILL
XFILL_72_DFFSR_236 gnd vdd FILL
XFILL_21_DFFSR_3 gnd vdd FILL
XFILL_69_DFFSR_80 gnd vdd FILL
XFILL_72_DFFSR_247 gnd vdd FILL
XFILL_26_NOR3X1_13 gnd vdd FILL
XFILL_69_DFFSR_91 gnd vdd FILL
XFILL_72_DFFSR_258 gnd vdd FILL
XFILL_72_DFFSR_269 gnd vdd FILL
XFILL_26_NOR3X1_24 gnd vdd FILL
XFILL_26_NOR3X1_35 gnd vdd FILL
XFILL_65_6_2 gnd vdd FILL
XFILL_26_NOR3X1_46 gnd vdd FILL
XFILL_76_DFFSR_202 gnd vdd FILL
XFILL_76_DFFSR_213 gnd vdd FILL
XFILL_59_DFFSR_1 gnd vdd FILL
XFILL_64_1_1 gnd vdd FILL
XFILL_76_DFFSR_224 gnd vdd FILL
XFILL_76_DFFSR_235 gnd vdd FILL
XFILL_76_DFFSR_246 gnd vdd FILL
XFILL_1_NOR3X1_7 gnd vdd FILL
XFILL_76_DFFSR_257 gnd vdd FILL
XFILL_76_DFFSR_268 gnd vdd FILL
XFILL_31_CLKBUF1_9 gnd vdd FILL
XFILL_11_DFFSR_190 gnd vdd FILL
XFILL_34_2 gnd vdd FILL
XFILL_38_DFFSR_90 gnd vdd FILL
XFILL_27_1 gnd vdd FILL
XFILL_35_CLKBUF1_8 gnd vdd FILL
XFILL_20_CLKBUF1_19 gnd vdd FILL
XFILL_43_DFFSR_7 gnd vdd FILL
XFILL_5_MUX2X1_190 gnd vdd FILL
XFILL_1_NOR2X1_108 gnd vdd FILL
XFILL_1_NOR2X1_119 gnd vdd FILL
XFILL_11_NAND2X1_12 gnd vdd FILL
XFILL_11_NAND2X1_23 gnd vdd FILL
XFILL_11_NAND2X1_34 gnd vdd FILL
XFILL_11_NAND2X1_45 gnd vdd FILL
XFILL_1_OAI21X1_4 gnd vdd FILL
XFILL_11_NAND2X1_56 gnd vdd FILL
XFILL_11_NAND2X1_67 gnd vdd FILL
XFILL_56_6_2 gnd vdd FILL
XFILL_9_OAI22X1_17 gnd vdd FILL
XFILL_11_NAND2X1_78 gnd vdd FILL
XFILL_9_OAI22X1_28 gnd vdd FILL
XFILL_11_NAND2X1_89 gnd vdd FILL
XFILL_9_OAI22X1_39 gnd vdd FILL
XFILL_55_1_1 gnd vdd FILL
XFILL_43_DFFSR_202 gnd vdd FILL
XFILL_43_DFFSR_213 gnd vdd FILL
XFILL_5_OAI21X1_3 gnd vdd FILL
XFILL_43_DFFSR_224 gnd vdd FILL
XFILL_43_DFFSR_235 gnd vdd FILL
XFILL_2_NOR2X1_50 gnd vdd FILL
XFILL_2_NOR2X1_61 gnd vdd FILL
XFILL_43_DFFSR_246 gnd vdd FILL
XFILL_8_NAND3X1_60 gnd vdd FILL
XFILL_43_DFFSR_257 gnd vdd FILL
XFILL_2_NOR2X1_72 gnd vdd FILL
XFILL_43_DFFSR_268 gnd vdd FILL
XFILL_8_NAND3X1_71 gnd vdd FILL
XNAND3X1_108 DFFSR_8/Q BUFX4_7/Y NOR3X1_9/Y gnd OAI21X1_19/C vdd NAND3X1
XFILL_2_NOR2X1_83 gnd vdd FILL
XNAND3X1_119 NOR2X1_82/Y NOR2X1_83/Y NOR3X1_31/Y gnd NOR2X1_84/A vdd NAND3X1
XFILL_70_DFFSR_102 gnd vdd FILL
XFILL_2_NOR2X1_94 gnd vdd FILL
XFILL_8_NAND3X1_82 gnd vdd FILL
XFILL_47_DFFSR_201 gnd vdd FILL
XFILL_8_NAND3X1_93 gnd vdd FILL
XFILL_70_DFFSR_113 gnd vdd FILL
XFILL_47_DFFSR_212 gnd vdd FILL
XFILL_5_BUFX4_6 gnd vdd FILL
XFILL_70_DFFSR_124 gnd vdd FILL
XFILL_9_OAI21X1_2 gnd vdd FILL
XFILL_47_DFFSR_223 gnd vdd FILL
XFILL_47_DFFSR_234 gnd vdd FILL
XFILL_70_DFFSR_135 gnd vdd FILL
XFILL_70_DFFSR_146 gnd vdd FILL
XFILL_47_DFFSR_245 gnd vdd FILL
XFILL_70_DFFSR_157 gnd vdd FILL
XFILL_6_NOR2X1_60 gnd vdd FILL
XFILL_6_NOR2X1_71 gnd vdd FILL
XFILL_70_DFFSR_168 gnd vdd FILL
XFILL_47_DFFSR_256 gnd vdd FILL
XFILL_47_DFFSR_267 gnd vdd FILL
XFILL_15_AND2X2_8 gnd vdd FILL
XFILL_6_NOR2X1_82 gnd vdd FILL
XFILL_70_DFFSR_179 gnd vdd FILL
XFILL_2_OAI21X1_19 gnd vdd FILL
XFILL_11_AOI22X1_10 gnd vdd FILL
XFILL_74_DFFSR_101 gnd vdd FILL
XFILL_6_NOR2X1_93 gnd vdd FILL
XFILL_74_DFFSR_112 gnd vdd FILL
XFILL_74_DFFSR_123 gnd vdd FILL
XFILL_74_DFFSR_134 gnd vdd FILL
XFILL_74_DFFSR_145 gnd vdd FILL
XFILL_15_AOI21X1_12 gnd vdd FILL
XFILL_74_DFFSR_156 gnd vdd FILL
XFILL_15_AOI21X1_23 gnd vdd FILL
XFILL_74_DFFSR_167 gnd vdd FILL
XFILL_15_AOI21X1_34 gnd vdd FILL
XFILL_74_DFFSR_178 gnd vdd FILL
XFILL_15_AOI21X1_45 gnd vdd FILL
XFILL_1_NAND2X1_40 gnd vdd FILL
XFILL_78_DFFSR_100 gnd vdd FILL
XFILL_74_DFFSR_189 gnd vdd FILL
XFILL_15_AOI21X1_56 gnd vdd FILL
XFILL_15_AOI21X1_67 gnd vdd FILL
XFILL_1_NAND2X1_51 gnd vdd FILL
XFILL_78_DFFSR_111 gnd vdd FILL
XFILL_15_AOI21X1_78 gnd vdd FILL
XFILL_1_NAND2X1_62 gnd vdd FILL
XFILL_78_DFFSR_122 gnd vdd FILL
XFILL_12_BUFX4_14 gnd vdd FILL
XFILL_78_DFFSR_133 gnd vdd FILL
XFILL_1_NAND2X1_73 gnd vdd FILL
XFILL_12_BUFX4_25 gnd vdd FILL
XFILL_1_NAND2X1_84 gnd vdd FILL
XFILL_12_BUFX4_36 gnd vdd FILL
XFILL_78_DFFSR_144 gnd vdd FILL
XFILL_1_NAND2X1_95 gnd vdd FILL
XFILL_78_DFFSR_155 gnd vdd FILL
XFILL_12_BUFX4_47 gnd vdd FILL
XFILL_78_DFFSR_166 gnd vdd FILL
XFILL_12_BUFX4_58 gnd vdd FILL
XFILL_78_DFFSR_177 gnd vdd FILL
XFILL_12_BUFX4_69 gnd vdd FILL
XFILL_1_BUFX2_2 gnd vdd FILL
XFILL_78_DFFSR_188 gnd vdd FILL
XFILL_78_DFFSR_199 gnd vdd FILL
XFILL_6_NAND3X1_130 gnd vdd FILL
XFILL_2_NAND2X1_5 gnd vdd FILL
XFILL_47_6_2 gnd vdd FILL
XFILL_60_DFFSR_1 gnd vdd FILL
XFILL_46_1_1 gnd vdd FILL
XFILL_6_INVX1_15 gnd vdd FILL
XFILL_6_NAND2X1_4 gnd vdd FILL
XFILL_10_DFFSR_202 gnd vdd FILL
XFILL_6_INVX1_26 gnd vdd FILL
XFILL_8_INVX8_4 gnd vdd FILL
XFILL_6_INVX1_37 gnd vdd FILL
XFILL_10_DFFSR_213 gnd vdd FILL
XFILL_18_MUX2X1_106 gnd vdd FILL
XFILL_18_MUX2X1_117 gnd vdd FILL
XFILL_6_INVX1_48 gnd vdd FILL
XFILL_7_AND2X2_7 gnd vdd FILL
XFILL_10_DFFSR_224 gnd vdd FILL
XFILL_10_DFFSR_235 gnd vdd FILL
XFILL_6_INVX1_59 gnd vdd FILL
XFILL_18_MUX2X1_128 gnd vdd FILL
XFILL_5_AOI21X1_40 gnd vdd FILL
XFILL_18_MUX2X1_139 gnd vdd FILL
XFILL_10_DFFSR_246 gnd vdd FILL
XFILL_2_MUX2X1_90 gnd vdd FILL
XFILL_5_AOI21X1_51 gnd vdd FILL
XFILL_10_DFFSR_257 gnd vdd FILL
XFILL_10_DFFSR_268 gnd vdd FILL
XFILL_15_OAI22X1_20 gnd vdd FILL
XFILL_5_AOI21X1_62 gnd vdd FILL
XFILL_5_AOI21X1_73 gnd vdd FILL
XFILL_15_OAI22X1_31 gnd vdd FILL
XFILL_14_DFFSR_201 gnd vdd FILL
XFILL_15_OAI22X1_42 gnd vdd FILL
XFILL_11_NAND3X1_1 gnd vdd FILL
XFILL_30_5_2 gnd vdd FILL
XFILL_14_DFFSR_212 gnd vdd FILL
XFILL_14_DFFSR_223 gnd vdd FILL
XFILL_14_DFFSR_234 gnd vdd FILL
XFILL_14_DFFSR_245 gnd vdd FILL
XFILL_25_DFFSR_4 gnd vdd FILL
XDFFSR_106 DFFSR_106/Q DFFSR_73/CLK DFFSR_73/R vdd DFFSR_106/D gnd vdd DFFSR
XFILL_8_NOR2X1_150 gnd vdd FILL
XFILL_14_DFFSR_256 gnd vdd FILL
XFILL_4_BUFX4_13 gnd vdd FILL
XFILL_8_NOR2X1_161 gnd vdd FILL
XFILL_14_DFFSR_267 gnd vdd FILL
XDFFSR_117 INVX1_179/A CLKBUF1_31/Y DFFSR_53/R vdd DFFSR_117/D gnd vdd DFFSR
XFILL_82_DFFSR_5 gnd vdd FILL
XFILL_4_BUFX4_24 gnd vdd FILL
XDFFSR_128 INVX1_172/A DFFSR_64/CLK DFFSR_64/R vdd DFFSR_128/D gnd vdd DFFSR
XFILL_8_NOR2X1_172 gnd vdd FILL
XFILL_41_DFFSR_101 gnd vdd FILL
XFILL_4_BUFX4_35 gnd vdd FILL
XFILL_8_NOR2X1_183 gnd vdd FILL
XDFFSR_139 DFFSR_139/Q DFFSR_55/CLK DFFSR_58/R vdd DFFSR_139/D gnd vdd DFFSR
XFILL_18_DFFSR_200 gnd vdd FILL
XFILL_4_BUFX4_46 gnd vdd FILL
XFILL_41_DFFSR_112 gnd vdd FILL
XFILL_18_DFFSR_211 gnd vdd FILL
XFILL_4_BUFX4_57 gnd vdd FILL
XFILL_8_NOR2X1_194 gnd vdd FILL
XFILL_18_DFFSR_222 gnd vdd FILL
XFILL_1_INVX2_2 gnd vdd FILL
XFILL_41_DFFSR_123 gnd vdd FILL
XFILL_41_DFFSR_134 gnd vdd FILL
XFILL_4_BUFX4_68 gnd vdd FILL
XFILL_18_DFFSR_233 gnd vdd FILL
XFILL_41_DFFSR_145 gnd vdd FILL
XFILL_18_DFFSR_244 gnd vdd FILL
XFILL_4_BUFX4_79 gnd vdd FILL
XFILL_41_DFFSR_156 gnd vdd FILL
XFILL_18_DFFSR_255 gnd vdd FILL
XFILL_41_DFFSR_167 gnd vdd FILL
XFILL_18_DFFSR_266 gnd vdd FILL
XFILL_41_DFFSR_178 gnd vdd FILL
XFILL_45_DFFSR_100 gnd vdd FILL
XFILL_41_DFFSR_189 gnd vdd FILL
XFILL_45_DFFSR_111 gnd vdd FILL
XFILL_45_DFFSR_122 gnd vdd FILL
XFILL_6_AOI21X1_9 gnd vdd FILL
XFILL_45_DFFSR_133 gnd vdd FILL
XFILL_45_DFFSR_144 gnd vdd FILL
XFILL_45_DFFSR_155 gnd vdd FILL
XFILL_45_DFFSR_166 gnd vdd FILL
XFILL_45_DFFSR_177 gnd vdd FILL
XFILL_45_DFFSR_188 gnd vdd FILL
XFILL_8_MUX2X1_101 gnd vdd FILL
XFILL_8_MUX2X1_112 gnd vdd FILL
XFILL_49_DFFSR_110 gnd vdd FILL
XFILL_45_DFFSR_199 gnd vdd FILL
XFILL_8_MUX2X1_123 gnd vdd FILL
XFILL_49_DFFSR_121 gnd vdd FILL
XFILL_49_DFFSR_132 gnd vdd FILL
XFILL_8_MUX2X1_134 gnd vdd FILL
XFILL_8_MUX2X1_145 gnd vdd FILL
XFILL_47_DFFSR_8 gnd vdd FILL
XFILL_49_DFFSR_143 gnd vdd FILL
XNOR3X1_17 NOR3X1_17/A NOR3X1_17/B NOR3X1_17/C gnd NOR3X1_17/Y vdd NOR3X1
XFILL_11_AND2X2_1 gnd vdd FILL
XFILL_49_DFFSR_154 gnd vdd FILL
XFILL_11_AOI22X1_6 gnd vdd FILL
XFILL_8_MUX2X1_156 gnd vdd FILL
XNOR3X1_28 NOR3X1_28/A NOR3X1_28/B NOR3X1_28/C gnd NOR3X1_28/Y vdd NOR3X1
XFILL_38_6_2 gnd vdd FILL
XFILL_49_DFFSR_165 gnd vdd FILL
XFILL_8_MUX2X1_167 gnd vdd FILL
XFILL_8_MUX2X1_178 gnd vdd FILL
XNOR3X1_39 INVX1_90/Y NOR3X1_49/B NOR3X1_39/C gnd NOR3X1_42/B vdd NOR3X1
XFILL_49_DFFSR_176 gnd vdd FILL
XFILL_8_MUX2X1_189 gnd vdd FILL
XFILL_49_DFFSR_187 gnd vdd FILL
XFILL_37_1_1 gnd vdd FILL
XFILL_49_DFFSR_198 gnd vdd FILL
XFILL_9_OAI21X1_50 gnd vdd FILL
XFILL_15_AOI22X1_5 gnd vdd FILL
XFILL_19_AOI22X1_4 gnd vdd FILL
XFILL_21_5_2 gnd vdd FILL
XFILL_20_0_1 gnd vdd FILL
XFILL_39_DFFSR_13 gnd vdd FILL
XFILL_39_DFFSR_24 gnd vdd FILL
XFILL_39_DFFSR_35 gnd vdd FILL
XFILL_39_DFFSR_46 gnd vdd FILL
XFILL_54_10 gnd vdd FILL
XFILL_39_DFFSR_57 gnd vdd FILL
XFILL_39_DFFSR_68 gnd vdd FILL
XFILL_39_DFFSR_79 gnd vdd FILL
XFILL_79_DFFSR_12 gnd vdd FILL
XFILL_79_DFFSR_23 gnd vdd FILL
XFILL_79_DFFSR_34 gnd vdd FILL
XFILL_79_DFFSR_45 gnd vdd FILL
XFILL_79_DFFSR_56 gnd vdd FILL
XFILL_10_NOR2X1_8 gnd vdd FILL
XFILL_79_DFFSR_67 gnd vdd FILL
XFILL_79_DFFSR_78 gnd vdd FILL
XFILL_79_DFFSR_89 gnd vdd FILL
XFILL_2_INVX1_30 gnd vdd FILL
XFILL_12_DFFSR_100 gnd vdd FILL
XFILL_12_DFFSR_111 gnd vdd FILL
XFILL_2_INVX1_41 gnd vdd FILL
XFILL_2_INVX1_52 gnd vdd FILL
XFILL_12_DFFSR_122 gnd vdd FILL
XFILL_9_BUFX4_7 gnd vdd FILL
XFILL_2_INVX1_63 gnd vdd FILL
XFILL_12_DFFSR_133 gnd vdd FILL
XFILL_2_INVX1_74 gnd vdd FILL
XFILL_12_DFFSR_144 gnd vdd FILL
XFILL_48_DFFSR_11 gnd vdd FILL
XFILL_2_INVX1_85 gnd vdd FILL
XFILL_12_DFFSR_155 gnd vdd FILL
XFILL_48_DFFSR_22 gnd vdd FILL
XFILL_2_INVX1_96 gnd vdd FILL
XFILL_12_DFFSR_166 gnd vdd FILL
XFILL_48_DFFSR_33 gnd vdd FILL
XFILL_19_NOR3X1_8 gnd vdd FILL
XFILL_48_DFFSR_44 gnd vdd FILL
XFILL_1_CLKBUF1_9 gnd vdd FILL
XFILL_12_DFFSR_177 gnd vdd FILL
XFILL_48_DFFSR_55 gnd vdd FILL
XFILL_12_DFFSR_188 gnd vdd FILL
XFILL_48_DFFSR_66 gnd vdd FILL
XFILL_16_DFFSR_110 gnd vdd FILL
XFILL_12_DFFSR_199 gnd vdd FILL
XFILL_48_DFFSR_77 gnd vdd FILL
XFILL_0_NAND3X1_15 gnd vdd FILL
XFILL_16_DFFSR_121 gnd vdd FILL
XFILL_29_6_2 gnd vdd FILL
XFILL_16_DFFSR_132 gnd vdd FILL
XFILL_4_6_2 gnd vdd FILL
XFILL_48_DFFSR_88 gnd vdd FILL
XFILL_48_DFFSR_99 gnd vdd FILL
XFILL_0_NAND3X1_26 gnd vdd FILL
XFILL_16_DFFSR_143 gnd vdd FILL
XFILL_0_NAND3X1_37 gnd vdd FILL
XFILL_28_1_1 gnd vdd FILL
XFILL_16_DFFSR_154 gnd vdd FILL
XFILL_3_1_1 gnd vdd FILL
XFILL_0_NAND3X1_48 gnd vdd FILL
XFILL_0_NAND3X1_59 gnd vdd FILL
XFILL_16_DFFSR_165 gnd vdd FILL
XFILL_16_DFFSR_176 gnd vdd FILL
XFILL_4_NAND2X1_17 gnd vdd FILL
XFILL_4_NAND2X1_28 gnd vdd FILL
XFILL_5_CLKBUF1_8 gnd vdd FILL
XFILL_17_DFFSR_10 gnd vdd FILL
XFILL_16_DFFSR_187 gnd vdd FILL
XFILL_0_BUFX4_50 gnd vdd FILL
XFILL_4_NAND2X1_39 gnd vdd FILL
XFILL_17_DFFSR_21 gnd vdd FILL
XFILL_16_DFFSR_198 gnd vdd FILL
XFILL_0_BUFX4_61 gnd vdd FILL
XFILL_0_BUFX4_72 gnd vdd FILL
XFILL_17_DFFSR_32 gnd vdd FILL
XFILL_17_DFFSR_43 gnd vdd FILL
XFILL_0_BUFX4_83 gnd vdd FILL
XFILL_17_DFFSR_54 gnd vdd FILL
XFILL_17_DFFSR_65 gnd vdd FILL
XFILL_0_BUFX4_94 gnd vdd FILL
XFILL_1_BUFX4_103 gnd vdd FILL
XFILL_17_DFFSR_76 gnd vdd FILL
XFILL_9_CLKBUF1_7 gnd vdd FILL
XFILL_17_DFFSR_87 gnd vdd FILL
XFILL_12_NOR3X1_11 gnd vdd FILL
XFILL_17_DFFSR_98 gnd vdd FILL
XFILL_5_BUFX2_3 gnd vdd FILL
XFILL_14_MUX2X1_170 gnd vdd FILL
XFILL_57_DFFSR_20 gnd vdd FILL
XFILL_12_NOR3X1_22 gnd vdd FILL
XFILL_12_NOR3X1_33 gnd vdd FILL
XFILL_14_MUX2X1_181 gnd vdd FILL
XFILL_12_NOR3X1_44 gnd vdd FILL
XFILL_12_5_2 gnd vdd FILL
XFILL_57_DFFSR_31 gnd vdd FILL
XFILL_62_DFFSR_200 gnd vdd FILL
XFILL_28_NOR3X1_6 gnd vdd FILL
XFILL_57_DFFSR_42 gnd vdd FILL
XFILL_14_MUX2X1_192 gnd vdd FILL
XFILL_62_DFFSR_211 gnd vdd FILL
XFILL_57_DFFSR_53 gnd vdd FILL
XFILL_62_DFFSR_222 gnd vdd FILL
XFILL_11_0_1 gnd vdd FILL
XFILL_57_DFFSR_64 gnd vdd FILL
XFILL_62_DFFSR_233 gnd vdd FILL
XFILL_5_BUFX4_102 gnd vdd FILL
XFILL_57_DFFSR_75 gnd vdd FILL
XFILL_62_DFFSR_244 gnd vdd FILL
XFILL_16_NOR3X1_10 gnd vdd FILL
XFILL_57_DFFSR_86 gnd vdd FILL
XFILL_62_DFFSR_255 gnd vdd FILL
XFILL_57_DFFSR_97 gnd vdd FILL
XFILL_62_DFFSR_266 gnd vdd FILL
XFILL_16_NOR3X1_21 gnd vdd FILL
XFILL_16_NOR3X1_32 gnd vdd FILL
XFILL_16_NOR3X1_43 gnd vdd FILL
XFILL_2_NOR2X1_7 gnd vdd FILL
XFILL_64_DFFSR_2 gnd vdd FILL
XFILL_66_DFFSR_210 gnd vdd FILL
XFILL_66_DFFSR_221 gnd vdd FILL
XFILL_9_BUFX4_101 gnd vdd FILL
XFILL_26_DFFSR_30 gnd vdd FILL
XFILL_66_DFFSR_232 gnd vdd FILL
XFILL_66_DFFSR_243 gnd vdd FILL
XFILL_26_DFFSR_41 gnd vdd FILL
XFILL_66_DFFSR_254 gnd vdd FILL
XFILL_26_DFFSR_52 gnd vdd FILL
XFILL_26_DFFSR_63 gnd vdd FILL
XFILL_66_DFFSR_265 gnd vdd FILL
XFILL_26_DFFSR_74 gnd vdd FILL
XFILL_21_CLKBUF1_6 gnd vdd FILL
XFILL_26_DFFSR_85 gnd vdd FILL
XFILL_26_DFFSR_96 gnd vdd FILL
XFILL_8_AOI21X1_17 gnd vdd FILL
XFILL_8_AOI21X1_28 gnd vdd FILL
XFILL_66_DFFSR_40 gnd vdd FILL
XFILL_8_AOI21X1_39 gnd vdd FILL
XFILL_1_MUX2X1_5 gnd vdd FILL
XFILL_66_DFFSR_51 gnd vdd FILL
XFILL_18_OAI22X1_19 gnd vdd FILL
XFILL_66_DFFSR_62 gnd vdd FILL
XFILL_25_CLKBUF1_5 gnd vdd FILL
XFILL_66_DFFSR_73 gnd vdd FILL
XFILL_66_DFFSR_84 gnd vdd FILL
XFILL_66_DFFSR_95 gnd vdd FILL
XFILL_3_NOR2X1_15 gnd vdd FILL
XFILL_3_NOR2X1_26 gnd vdd FILL
XNAND3X1_50 AOI22X1_4/Y NAND3X1_50/B NOR3X1_50/Y gnd NOR3X1_3/A vdd NAND3X1
XFILL_3_NOR2X1_37 gnd vdd FILL
XNAND3X1_61 BUFX4_57/Y AND2X2_5/B NOR2X1_42/Y gnd OAI22X1_6/D vdd NAND3X1
XFILL_9_DFFSR_20 gnd vdd FILL
XFILL_3_NOR2X1_48 gnd vdd FILL
XFILL_29_DFFSR_5 gnd vdd FILL
XFILL_3_NOR2X1_59 gnd vdd FILL
XFILL_9_DFFSR_31 gnd vdd FILL
XNAND3X1_72 AND2X2_6/A AND2X2_5/B BUFX4_103/Y gnd OAI22X1_5/D vdd NAND3X1
XFILL_86_DFFSR_6 gnd vdd FILL
XFILL_29_CLKBUF1_4 gnd vdd FILL
XNAND3X1_83 DFFSR_29/Q NAND3X1_7/B NOR2X1_37/Y gnd OAI21X1_8/C vdd NAND3X1
XFILL_9_DFFSR_42 gnd vdd FILL
XFILL_7_NAND3X1_120 gnd vdd FILL
XNAND3X1_94 DFFSR_82/Q BUFX4_1/Y NOR2X1_44/Y gnd OAI21X1_15/C vdd NAND3X1
XFILL_7_NAND3X1_131 gnd vdd FILL
XFILL_9_DFFSR_53 gnd vdd FILL
XFILL_19_1_1 gnd vdd FILL
XFILL_9_DFFSR_64 gnd vdd FILL
XFILL_9_DFFSR_75 gnd vdd FILL
XFILL_7_NOR2X1_14 gnd vdd FILL
XFILL_35_DFFSR_50 gnd vdd FILL
XFILL_9_DFFSR_86 gnd vdd FILL
XFILL_7_NOR2X1_25 gnd vdd FILL
XFILL_5_INVX2_3 gnd vdd FILL
XFILL_7_NOR2X1_36 gnd vdd FILL
XNOR2X1_50 NOR3X1_29/B NOR3X1_6/C gnd NOR2X1_50/Y vdd NOR2X1
XFILL_35_DFFSR_61 gnd vdd FILL
XFILL_35_DFFSR_72 gnd vdd FILL
XFILL_9_DFFSR_97 gnd vdd FILL
XFILL_35_DFFSR_83 gnd vdd FILL
XFILL_7_NOR2X1_47 gnd vdd FILL
XNOR2X1_61 OAI21X1_8/Y NOR2X1_61/B gnd NOR2X1_61/Y vdd NOR2X1
XFILL_7_NOR2X1_58 gnd vdd FILL
XFILL_35_DFFSR_94 gnd vdd FILL
XFILL_11_OAI22X1_9 gnd vdd FILL
XNOR2X1_72 INVX1_73/Y OAI22X1_1/B gnd NOR3X1_25/B vdd NOR2X1
XFILL_62_4_2 gnd vdd FILL
XFILL_7_NOR2X1_69 gnd vdd FILL
XNOR2X1_83 NOR2X1_83/A NOR2X1_83/B gnd NOR2X1_83/Y vdd NOR2X1
XNOR2X1_94 NOR2X1_94/A NOR2X1_94/B gnd NOR2X1_94/Y vdd NOR2X1
XFILL_0_NOR2X1_105 gnd vdd FILL
XFILL_0_NOR2X1_116 gnd vdd FILL
XFILL_75_DFFSR_60 gnd vdd FILL
XFILL_0_NOR2X1_127 gnd vdd FILL
XFILL_75_DFFSR_71 gnd vdd FILL
XFILL_75_DFFSR_82 gnd vdd FILL
XFILL_0_NOR2X1_138 gnd vdd FILL
XFILL_0_NOR2X1_149 gnd vdd FILL
XFILL_15_OAI22X1_8 gnd vdd FILL
XFILL_75_DFFSR_93 gnd vdd FILL
XFILL_3_INVX1_1 gnd vdd FILL
XFILL_11_4 gnd vdd FILL
XFILL_10_NAND2X1_20 gnd vdd FILL
XFILL_79_DFFSR_109 gnd vdd FILL
XFILL_10_NAND2X1_31 gnd vdd FILL
XFILL_10_NAND2X1_42 gnd vdd FILL
XFILL_10_NAND2X1_53 gnd vdd FILL
XFILL_15_NOR3X1_1 gnd vdd FILL
XFILL_10_NAND2X1_64 gnd vdd FILL
XFILL_19_OAI22X1_7 gnd vdd FILL
XFILL_8_OAI22X1_14 gnd vdd FILL
XFILL_10_NAND2X1_75 gnd vdd FILL
XFILL_8_OAI22X1_25 gnd vdd FILL
XFILL_44_DFFSR_70 gnd vdd FILL
XFILL_8_OAI22X1_36 gnd vdd FILL
XFILL_10_NAND2X1_86 gnd vdd FILL
XFILL_8_OAI22X1_47 gnd vdd FILL
XFILL_44_DFFSR_81 gnd vdd FILL
XFILL_44_DFFSR_92 gnd vdd FILL
XFILL_33_DFFSR_210 gnd vdd FILL
XFILL_33_DFFSR_221 gnd vdd FILL
XFILL_33_DFFSR_232 gnd vdd FILL
XFILL_33_DFFSR_243 gnd vdd FILL
XFILL_33_DFFSR_254 gnd vdd FILL
XFILL_84_DFFSR_80 gnd vdd FILL
XFILL_33_DFFSR_265 gnd vdd FILL
XFILL_84_DFFSR_91 gnd vdd FILL
XFILL_60_DFFSR_110 gnd vdd FILL
XFILL_7_NAND3X1_90 gnd vdd FILL
XFILL_60_DFFSR_121 gnd vdd FILL
XFILL_13_DFFSR_80 gnd vdd FILL
XFILL_5_NOR2X1_205 gnd vdd FILL
XFILL_37_DFFSR_220 gnd vdd FILL
XFILL_60_DFFSR_132 gnd vdd FILL
XFILL_37_DFFSR_231 gnd vdd FILL
XFILL_60_DFFSR_143 gnd vdd FILL
XFILL_37_DFFSR_242 gnd vdd FILL
XFILL_13_DFFSR_91 gnd vdd FILL
XFILL_60_DFFSR_154 gnd vdd FILL
XFILL_37_DFFSR_253 gnd vdd FILL
XFILL_60_DFFSR_165 gnd vdd FILL
XNAND2X1_5 AND2X2_8/B INVX2_1/A gnd NAND2X1_5/Y vdd NAND2X1
XFILL_37_DFFSR_264 gnd vdd FILL
XFILL_3_MUX2X1_11 gnd vdd FILL
XFILL_60_DFFSR_176 gnd vdd FILL
XFILL_37_DFFSR_275 gnd vdd FILL
XFILL_3_MUX2X1_22 gnd vdd FILL
XFILL_1_OAI21X1_16 gnd vdd FILL
XFILL_60_DFFSR_187 gnd vdd FILL
XFILL_3_MUX2X1_33 gnd vdd FILL
XFILL_19_CLKBUF1_12 gnd vdd FILL
XFILL_1_OAI21X1_27 gnd vdd FILL
XFILL_60_DFFSR_198 gnd vdd FILL
XFILL_64_DFFSR_120 gnd vdd FILL
XFILL_19_CLKBUF1_23 gnd vdd FILL
XFILL_1_OAI21X1_38 gnd vdd FILL
XFILL_3_MUX2X1_44 gnd vdd FILL
XFILL_64_DFFSR_131 gnd vdd FILL
XFILL_19_CLKBUF1_34 gnd vdd FILL
XFILL_1_OAI21X1_49 gnd vdd FILL
XFILL_3_MUX2X1_55 gnd vdd FILL
XFILL_53_DFFSR_90 gnd vdd FILL
XFILL_3_MUX2X1_66 gnd vdd FILL
XFILL_3_MUX2X1_77 gnd vdd FILL
XFILL_64_DFFSR_142 gnd vdd FILL
XFILL_14_AOI21X1_20 gnd vdd FILL
XFILL_64_DFFSR_153 gnd vdd FILL
XFILL_3_MUX2X1_88 gnd vdd FILL
XFILL_14_AOI21X1_31 gnd vdd FILL
XFILL_64_DFFSR_164 gnd vdd FILL
XFILL_3_MUX2X1_99 gnd vdd FILL
XFILL_64_DFFSR_175 gnd vdd FILL
XFILL_7_MUX2X1_10 gnd vdd FILL
XFILL_7_MUX2X1_21 gnd vdd FILL
XFILL_14_AOI21X1_42 gnd vdd FILL
XFILL_64_DFFSR_186 gnd vdd FILL
XFILL_7_MUX2X1_32 gnd vdd FILL
XFILL_14_AOI21X1_53 gnd vdd FILL
XFILL_64_DFFSR_197 gnd vdd FILL
XFILL_14_AOI21X1_64 gnd vdd FILL
XFILL_7_MUX2X1_43 gnd vdd FILL
XFILL_53_4_2 gnd vdd FILL
XFILL_14_AOI21X1_75 gnd vdd FILL
XFILL_68_DFFSR_130 gnd vdd FILL
XFILL_7_MUX2X1_54 gnd vdd FILL
XFILL_0_NAND2X1_70 gnd vdd FILL
XFILL_0_NAND2X1_81 gnd vdd FILL
XNOR2X1_140 BUFX2_8/A INVX1_140/Y gnd NAND3X1_1/B vdd NOR2X1
XFILL_7_MUX2X1_65 gnd vdd FILL
XFILL_68_DFFSR_141 gnd vdd FILL
XMUX2X1_90 MUX2X1_1/A MUX2X1_90/B NOR2X1_57/Y gnd MUX2X1_90/Y vdd MUX2X1
XFILL_7_MUX2X1_76 gnd vdd FILL
XNOR2X1_151 DFFSR_100/Q NOR2X1_153/B gnd NOR2X1_151/Y vdd NOR2X1
XFILL_0_NAND2X1_92 gnd vdd FILL
XFILL_68_DFFSR_152 gnd vdd FILL
XFILL_7_MUX2X1_87 gnd vdd FILL
XNOR2X1_162 OR2X2_1/B NAND2X1_3/Y gnd NOR2X1_162/Y vdd NOR2X1
XNOR2X1_173 DFFSR_40/Q MUX2X1_9/S gnd NOR2X1_173/Y vdd NOR2X1
XFILL_68_DFFSR_163 gnd vdd FILL
XFILL_68_DFFSR_174 gnd vdd FILL
XFILL_7_MUX2X1_98 gnd vdd FILL
XNOR2X1_184 DFFSR_26/Q MUX2X1_16/S gnd NOR2X1_184/Y vdd NOR2X1
XFILL_68_DFFSR_185 gnd vdd FILL
XNOR2X1_195 DFFSR_18/Q NOR2X1_195/B gnd NOR2X1_195/Y vdd NOR2X1
XFILL_68_DFFSR_196 gnd vdd FILL
XFILL_19_DFFSR_209 gnd vdd FILL
XFILL_46_DFFSR_109 gnd vdd FILL
XMUX2X1_102 NOR3X1_26/A BUFX4_68/Y NAND2X1_16/Y gnd DFFSR_24/D vdd MUX2X1
XMUX2X1_113 BUFX4_80/Y OAI21X1_3/A NOR2X1_128/Y gnd DFFSR_143/D vdd MUX2X1
XMUX2X1_124 BUFX4_76/Y INVX1_168/Y NOR2X1_136/Y gnd DFFSR_132/D vdd MUX2X1
XFILL_5_DFFSR_90 gnd vdd FILL
XMUX2X1_135 BUFX4_87/Y INVX1_179/Y NOR2X1_139/Y gnd DFFSR_117/D vdd MUX2X1
XFILL_23_MUX2X1_30 gnd vdd FILL
XFILL_9_CLKBUF1_40 gnd vdd FILL
XFILL_17_MUX2X1_103 gnd vdd FILL
XMUX2X1_146 BUFX4_74/Y INVX1_190/Y NOR2X1_142/Y gnd DFFSR_109/D vdd MUX2X1
XFILL_17_MUX2X1_114 gnd vdd FILL
XFILL_23_MUX2X1_41 gnd vdd FILL
XMUX2X1_157 BUFX4_81/Y INVX1_201/Y NOR2X1_156/Y gnd DFFSR_85/D vdd MUX2X1
XFILL_17_MUX2X1_125 gnd vdd FILL
XFILL_23_MUX2X1_52 gnd vdd FILL
XMUX2X1_168 BUFX4_74/Y INVX1_213/Y NOR2X1_164/Y gnd DFFSR_74/D vdd MUX2X1
XFILL_17_MUX2X1_136 gnd vdd FILL
XFILL_23_MUX2X1_63 gnd vdd FILL
XMUX2X1_179 BUFX4_87/Y INVX1_224/Y NOR2X1_167/Y gnd DFFSR_59/D vdd MUX2X1
XFILL_23_MUX2X1_74 gnd vdd FILL
XFILL_23_MUX2X1_85 gnd vdd FILL
XFILL_17_MUX2X1_147 gnd vdd FILL
XFILL_17_MUX2X1_158 gnd vdd FILL
XFILL_4_AOI21X1_70 gnd vdd FILL
XFILL_23_MUX2X1_96 gnd vdd FILL
XFILL_9_BUFX2_4 gnd vdd FILL
XFILL_17_MUX2X1_169 gnd vdd FILL
XFILL_4_AOI21X1_81 gnd vdd FILL
XINVX1_20 INVX1_20/A gnd MUX2X1_7/A vdd INVX1
XFILL_14_OAI22X1_50 gnd vdd FILL
XINVX1_31 INVX1_31/A gnd INVX1_31/Y vdd INVX1
XINVX1_42 INVX1_42/A gnd INVX1_42/Y vdd INVX1
XINVX1_53 INVX1_53/A gnd INVX1_53/Y vdd INVX1
XFILL_30_DFFSR_5 gnd vdd FILL
XINVX1_64 INVX1_64/A gnd INVX1_64/Y vdd INVX1
XINVX1_75 INVX1_75/A gnd INVX1_75/Y vdd INVX1
XINVX1_86 INVX1_86/A gnd INVX1_86/Y vdd INVX1
XINVX1_97 INVX1_97/A gnd INVX1_97/Y vdd INVX1
XFILL_7_NOR2X1_180 gnd vdd FILL
XFILL_68_DFFSR_3 gnd vdd FILL
XFILL_7_NOR2X1_191 gnd vdd FILL
XFILL_31_DFFSR_120 gnd vdd FILL
XFILL_31_DFFSR_131 gnd vdd FILL
XFILL_3_INVX1_19 gnd vdd FILL
XFILL_31_DFFSR_142 gnd vdd FILL
XFILL_31_DFFSR_153 gnd vdd FILL
XFILL_44_4_2 gnd vdd FILL
XFILL_31_DFFSR_164 gnd vdd FILL
XFILL_31_DFFSR_175 gnd vdd FILL
XFILL_31_DFFSR_186 gnd vdd FILL
XFILL_31_DFFSR_197 gnd vdd FILL
XFILL_35_DFFSR_130 gnd vdd FILL
XFILL_35_DFFSR_141 gnd vdd FILL
XFILL_35_DFFSR_152 gnd vdd FILL
XFILL_35_DFFSR_163 gnd vdd FILL
XFILL_35_DFFSR_174 gnd vdd FILL
XFILL_35_DFFSR_185 gnd vdd FILL
XFILL_35_DFFSR_196 gnd vdd FILL
XFILL_7_MUX2X1_120 gnd vdd FILL
XFILL_1_BUFX4_17 gnd vdd FILL
XFILL_52_DFFSR_9 gnd vdd FILL
XFILL_1_BUFX4_28 gnd vdd FILL
XFILL_7_MUX2X1_131 gnd vdd FILL
XFILL_39_DFFSR_140 gnd vdd FILL
XFILL_7_MUX2X1_142 gnd vdd FILL
XFILL_1_BUFX4_39 gnd vdd FILL
XFILL_7_MUX2X1_153 gnd vdd FILL
XFILL_39_DFFSR_151 gnd vdd FILL
XFILL_39_DFFSR_162 gnd vdd FILL
XFILL_7_MUX2X1_164 gnd vdd FILL
XFILL_7_MUX2X1_175 gnd vdd FILL
XFILL_39_DFFSR_173 gnd vdd FILL
XFILL_39_DFFSR_184 gnd vdd FILL
XFILL_7_MUX2X1_186 gnd vdd FILL
XFILL_39_DFFSR_195 gnd vdd FILL
XFILL_31_NOR3X1_20 gnd vdd FILL
XFILL_13_DFFSR_109 gnd vdd FILL
XFILL_31_NOR3X1_31 gnd vdd FILL
XFILL_31_NOR3X1_42 gnd vdd FILL
XFILL_81_DFFSR_220 gnd vdd FILL
XNOR2X1_8 NOR2X1_8/A NOR2X1_9/B gnd NOR2X1_8/Y vdd NOR2X1
XFILL_81_DFFSR_231 gnd vdd FILL
XFILL_81_DFFSR_242 gnd vdd FILL
XFILL_81_DFFSR_253 gnd vdd FILL
XFILL_81_DFFSR_264 gnd vdd FILL
XFILL_81_DFFSR_275 gnd vdd FILL
XFILL_17_DFFSR_108 gnd vdd FILL
XFILL_17_DFFSR_119 gnd vdd FILL
XFILL_7_INVX1_2 gnd vdd FILL
XFILL_85_DFFSR_230 gnd vdd FILL
XFILL_12_AOI21X1_4 gnd vdd FILL
XFILL_85_DFFSR_241 gnd vdd FILL
XFILL_85_DFFSR_252 gnd vdd FILL
XFILL_27_DFFSR_19 gnd vdd FILL
XFILL_85_DFFSR_263 gnd vdd FILL
XFILL_85_DFFSR_274 gnd vdd FILL
XFILL_66_5 gnd vdd FILL
XFILL_59_4 gnd vdd FILL
XFILL_1_INVX1_180 gnd vdd FILL
XFILL_8_NAND3X1_110 gnd vdd FILL
XFILL_8_NAND3X1_121 gnd vdd FILL
XFILL_67_DFFSR_18 gnd vdd FILL
XFILL_1_INVX1_191 gnd vdd FILL
XFILL_8_NAND3X1_132 gnd vdd FILL
XFILL_67_DFFSR_29 gnd vdd FILL
XFILL_63_7_0 gnd vdd FILL
XFILL_35_4_2 gnd vdd FILL
XFILL_63_DFFSR_209 gnd vdd FILL
XFILL_5_INVX1_190 gnd vdd FILL
XFILL_17_NOR3X1_19 gnd vdd FILL
XFILL_67_DFFSR_208 gnd vdd FILL
XFILL_67_DFFSR_219 gnd vdd FILL
XFILL_36_DFFSR_17 gnd vdd FILL
XFILL_36_DFFSR_28 gnd vdd FILL
XFILL_36_DFFSR_39 gnd vdd FILL
XAOI21X1_18 BUFX4_68/Y NOR2X1_161/B NOR2X1_159/Y gnd DFFSR_82/D vdd AOI21X1
XAOI21X1_29 MUX2X1_6/B MUX2X1_16/S NOR2X1_184/Y gnd DFFSR_26/D vdd AOI21X1
XFILL_76_DFFSR_16 gnd vdd FILL
XFILL_76_DFFSR_27 gnd vdd FILL
XFILL_76_DFFSR_38 gnd vdd FILL
XFILL_76_DFFSR_49 gnd vdd FILL
XFILL_3_NAND2X1_14 gnd vdd FILL
XFILL_19_MUX2X1_6 gnd vdd FILL
XFILL_3_NAND2X1_25 gnd vdd FILL
XFILL_3_NAND2X1_36 gnd vdd FILL
XFILL_3_NAND2X1_47 gnd vdd FILL
XFILL_3_NAND2X1_58 gnd vdd FILL
XFILL_3_NAND2X1_69 gnd vdd FILL
XFILL_0_AND2X2_4 gnd vdd FILL
XFILL_45_DFFSR_15 gnd vdd FILL
XFILL_45_DFFSR_26 gnd vdd FILL
XFILL_45_DFFSR_37 gnd vdd FILL
XFILL_45_DFFSR_48 gnd vdd FILL
XFILL_45_DFFSR_59 gnd vdd FILL
XFILL_52_DFFSR_230 gnd vdd FILL
XFILL_52_DFFSR_241 gnd vdd FILL
XFILL_85_DFFSR_14 gnd vdd FILL
XFILL_52_DFFSR_252 gnd vdd FILL
XFILL_85_DFFSR_25 gnd vdd FILL
XFILL_12_DFFSR_2 gnd vdd FILL
XFILL_52_DFFSR_263 gnd vdd FILL
XFILL_52_DFFSR_274 gnd vdd FILL
XFILL_85_DFFSR_36 gnd vdd FILL
XFILL_85_DFFSR_47 gnd vdd FILL
XFILL_85_DFFSR_58 gnd vdd FILL
XFILL_14_DFFSR_14 gnd vdd FILL
XFILL_29_CLKBUF1_13 gnd vdd FILL
XFILL_29_CLKBUF1_24 gnd vdd FILL
XFILL_85_DFFSR_69 gnd vdd FILL
XFILL_14_DFFSR_25 gnd vdd FILL
XFILL_29_CLKBUF1_35 gnd vdd FILL
XFILL_14_DFFSR_36 gnd vdd FILL
XFILL_56_DFFSR_240 gnd vdd FILL
XFILL_14_DFFSR_47 gnd vdd FILL
XFILL_54_7_0 gnd vdd FILL
XFILL_14_DFFSR_58 gnd vdd FILL
XFILL_56_DFFSR_251 gnd vdd FILL
XFILL_14_DFFSR_69 gnd vdd FILL
XFILL_26_4_2 gnd vdd FILL
XFILL_11_CLKBUF1_3 gnd vdd FILL
XFILL_56_DFFSR_262 gnd vdd FILL
XFILL_1_4_2 gnd vdd FILL
XFILL_56_DFFSR_273 gnd vdd FILL
XFILL_54_DFFSR_13 gnd vdd FILL
XFILL_54_DFFSR_24 gnd vdd FILL
XFILL_30_DFFSR_209 gnd vdd FILL
XFILL_7_AOI21X1_14 gnd vdd FILL
XOAI22X1_15 INVX1_55/Y OAI22X1_33/B INVX1_60/Y OAI22X1_33/D gnd NOR2X1_73/B vdd OAI22X1
XFILL_54_DFFSR_35 gnd vdd FILL
XFILL_7_AOI21X1_25 gnd vdd FILL
XOAI22X1_26 INVX1_23/Y NOR2X1_66/B INVX1_27/Y OAI22X1_26/D gnd NOR2X1_85/A vdd OAI22X1
XFILL_83_DFFSR_140 gnd vdd FILL
XFILL_54_DFFSR_46 gnd vdd FILL
XFILL_7_AOI21X1_36 gnd vdd FILL
XOAI22X1_37 INVX1_223/Y OAI22X1_9/B INVX1_227/Y OAI22X1_9/D gnd NOR2X1_99/B vdd OAI22X1
XFILL_54_DFFSR_57 gnd vdd FILL
XFILL_83_DFFSR_151 gnd vdd FILL
XFILL_7_AOI21X1_47 gnd vdd FILL
XFILL_83_DFFSR_162 gnd vdd FILL
XFILL_54_DFFSR_68 gnd vdd FILL
XOAI22X1_48 INVX1_211/Y OAI22X1_48/B INVX1_215/Y OAI22X1_48/D gnd NOR2X1_48/A vdd
+ OAI22X1
XFILL_83_DFFSR_173 gnd vdd FILL
XFILL_54_DFFSR_79 gnd vdd FILL
XFILL_17_OAI22X1_16 gnd vdd FILL
XFILL_7_AOI21X1_58 gnd vdd FILL
XFILL_15_CLKBUF1_2 gnd vdd FILL
XFILL_83_DFFSR_184 gnd vdd FILL
XFILL_7_AOI21X1_69 gnd vdd FILL
XFILL_17_OAI22X1_27 gnd vdd FILL
XFILL_3_DFFSR_210 gnd vdd FILL
XFILL_83_DFFSR_195 gnd vdd FILL
XFILL_17_OAI22X1_38 gnd vdd FILL
XFILL_34_DFFSR_208 gnd vdd FILL
XFILL_3_DFFSR_221 gnd vdd FILL
XFILL_17_OAI22X1_49 gnd vdd FILL
XFILL_34_DFFSR_219 gnd vdd FILL
XFILL_3_DFFSR_232 gnd vdd FILL
XFILL_3_DFFSR_243 gnd vdd FILL
XFILL_34_DFFSR_6 gnd vdd FILL
XFILL_23_DFFSR_12 gnd vdd FILL
XFILL_3_DFFSR_254 gnd vdd FILL
XFILL_87_DFFSR_150 gnd vdd FILL
XFILL_87_DFFSR_161 gnd vdd FILL
XFILL_23_DFFSR_23 gnd vdd FILL
XFILL_3_DFFSR_265 gnd vdd FILL
XFILL_19_CLKBUF1_1 gnd vdd FILL
XFILL_87_DFFSR_172 gnd vdd FILL
XFILL_23_DFFSR_34 gnd vdd FILL
XFILL_1_CLKBUF1_17 gnd vdd FILL
XFILL_1_CLKBUF1_28 gnd vdd FILL
XFILL_87_DFFSR_183 gnd vdd FILL
XFILL_87_DFFSR_194 gnd vdd FILL
XFILL_23_DFFSR_45 gnd vdd FILL
XFILL_1_CLKBUF1_39 gnd vdd FILL
XFILL_38_DFFSR_207 gnd vdd FILL
XFILL_23_DFFSR_56 gnd vdd FILL
XFILL_61_DFFSR_108 gnd vdd FILL
XFILL_23_DFFSR_67 gnd vdd FILL
XFILL_7_DFFSR_220 gnd vdd FILL
XFILL_61_DFFSR_119 gnd vdd FILL
XFILL_23_DFFSR_78 gnd vdd FILL
XFILL_38_DFFSR_218 gnd vdd FILL
XFILL_7_DFFSR_231 gnd vdd FILL
XFILL_23_DFFSR_89 gnd vdd FILL
XFILL_7_DFFSR_242 gnd vdd FILL
XFILL_38_DFFSR_229 gnd vdd FILL
XFILL_7_DFFSR_253 gnd vdd FILL
XFILL_63_DFFSR_11 gnd vdd FILL
XFILL_63_DFFSR_22 gnd vdd FILL
XFILL_7_DFFSR_264 gnd vdd FILL
XFILL_7_DFFSR_275 gnd vdd FILL
XFILL_63_DFFSR_33 gnd vdd FILL
XFILL_63_DFFSR_44 gnd vdd FILL
XFILL_65_DFFSR_107 gnd vdd FILL
XFILL_63_DFFSR_55 gnd vdd FILL
XFILL_63_DFFSR_66 gnd vdd FILL
XFILL_65_DFFSR_118 gnd vdd FILL
XFILL_63_DFFSR_77 gnd vdd FILL
XFILL_10_OAI21X1_18 gnd vdd FILL
XFILL_65_DFFSR_129 gnd vdd FILL
XFILL_10_OAI21X1_29 gnd vdd FILL
XFILL_9_5_2 gnd vdd FILL
XFILL_63_DFFSR_88 gnd vdd FILL
XFILL_63_DFFSR_99 gnd vdd FILL
XFILL_8_0_1 gnd vdd FILL
XFILL_6_DFFSR_13 gnd vdd FILL
XFILL_6_DFFSR_24 gnd vdd FILL
XFILL_8_MUX2X1_19 gnd vdd FILL
XFILL_6_DFFSR_35 gnd vdd FILL
XFILL_69_DFFSR_106 gnd vdd FILL
XFILL_32_DFFSR_10 gnd vdd FILL
XFILL_32_DFFSR_21 gnd vdd FILL
XFILL_6_DFFSR_46 gnd vdd FILL
XFILL_69_DFFSR_117 gnd vdd FILL
XFILL_6_DFFSR_57 gnd vdd FILL
XFILL_32_DFFSR_32 gnd vdd FILL
XFILL_69_DFFSR_128 gnd vdd FILL
XFILL_32_DFFSR_43 gnd vdd FILL
XFILL_6_DFFSR_68 gnd vdd FILL
XFILL_69_DFFSR_139 gnd vdd FILL
XFILL_6_DFFSR_79 gnd vdd FILL
XFILL_32_DFFSR_54 gnd vdd FILL
XFILL_0_AOI22X1_4 gnd vdd FILL
XFILL_12_OAI21X1_7 gnd vdd FILL
XFILL_7_OAI22X1_11 gnd vdd FILL
XFILL_32_DFFSR_65 gnd vdd FILL
XFILL_7_OAI22X1_22 gnd vdd FILL
XFILL_32_DFFSR_76 gnd vdd FILL
XFILL_7_OAI22X1_33 gnd vdd FILL
XFILL_7_OAI22X1_44 gnd vdd FILL
XFILL_32_DFFSR_87 gnd vdd FILL
XFILL_32_DFFSR_98 gnd vdd FILL
XFILL_0_INVX1_203 gnd vdd FILL
XFILL_45_7_0 gnd vdd FILL
XFILL_72_DFFSR_20 gnd vdd FILL
XFILL_0_INVX1_214 gnd vdd FILL
XFILL_72_DFFSR_31 gnd vdd FILL
XFILL_0_INVX1_225 gnd vdd FILL
XFILL_17_4_2 gnd vdd FILL
XFILL_72_DFFSR_42 gnd vdd FILL
XFILL_72_DFFSR_53 gnd vdd FILL
XFILL_4_AOI22X1_3 gnd vdd FILL
XFILL_23_DFFSR_240 gnd vdd FILL
XFILL_72_DFFSR_64 gnd vdd FILL
XFILL_23_DFFSR_251 gnd vdd FILL
XFILL_72_DFFSR_75 gnd vdd FILL
XFILL_72_DFFSR_86 gnd vdd FILL
XFILL_23_DFFSR_262 gnd vdd FILL
XFILL_4_INVX1_202 gnd vdd FILL
XFILL_23_DFFSR_273 gnd vdd FILL
XFILL_72_DFFSR_97 gnd vdd FILL
XFILL_20_MUX2X1_18 gnd vdd FILL
XFILL_20_MUX2X1_29 gnd vdd FILL
XFILL_4_INVX1_213 gnd vdd FILL
XFILL_4_NOR2X1_202 gnd vdd FILL
XFILL_4_INVX1_224 gnd vdd FILL
XFILL_8_AOI22X1_2 gnd vdd FILL
XFILL_50_DFFSR_140 gnd vdd FILL
XFILL_50_DFFSR_151 gnd vdd FILL
XFILL_27_DFFSR_250 gnd vdd FILL
XFILL_50_DFFSR_162 gnd vdd FILL
XFILL_41_DFFSR_30 gnd vdd FILL
XFILL_27_DFFSR_261 gnd vdd FILL
XFILL_50_DFFSR_173 gnd vdd FILL
XFILL_41_DFFSR_41 gnd vdd FILL
XFILL_12_NOR3X1_5 gnd vdd FILL
XFILL_50_DFFSR_184 gnd vdd FILL
XFILL_0_OAI21X1_13 gnd vdd FILL
XFILL_27_DFFSR_272 gnd vdd FILL
XFILL_41_DFFSR_52 gnd vdd FILL
XFILL_41_DFFSR_63 gnd vdd FILL
XFILL_0_OAI21X1_24 gnd vdd FILL
XFILL_50_DFFSR_195 gnd vdd FILL
XFILL_41_DFFSR_74 gnd vdd FILL
XFILL_18_CLKBUF1_20 gnd vdd FILL
XFILL_0_OAI21X1_35 gnd vdd FILL
XFILL_41_DFFSR_85 gnd vdd FILL
XFILL_18_CLKBUF1_31 gnd vdd FILL
XFILL_0_OAI21X1_46 gnd vdd FILL
XFILL_41_DFFSR_96 gnd vdd FILL
XFILL_18_CLKBUF1_42 gnd vdd FILL
XFILL_54_DFFSR_150 gnd vdd FILL
XFILL_54_DFFSR_161 gnd vdd FILL
XFILL_81_DFFSR_40 gnd vdd FILL
XFILL_54_DFFSR_172 gnd vdd FILL
XFILL_81_DFFSR_51 gnd vdd FILL
XFILL_54_DFFSR_183 gnd vdd FILL
XFILL_13_AOI21X1_50 gnd vdd FILL
XFILL_81_DFFSR_62 gnd vdd FILL
XFILL_81_DFFSR_73 gnd vdd FILL
XFILL_54_DFFSR_194 gnd vdd FILL
XFILL_13_AOI21X1_61 gnd vdd FILL
XFILL_81_DFFSR_84 gnd vdd FILL
XFILL_10_DFFSR_40 gnd vdd FILL
XFILL_13_AOI21X1_72 gnd vdd FILL
XFILL_81_DFFSR_95 gnd vdd FILL
XFILL_10_DFFSR_51 gnd vdd FILL
XFILL_10_DFFSR_62 gnd vdd FILL
XFILL_10_DFFSR_73 gnd vdd FILL
XFILL_58_DFFSR_160 gnd vdd FILL
XFILL_10_DFFSR_84 gnd vdd FILL
XFILL_58_DFFSR_171 gnd vdd FILL
XFILL_10_DFFSR_95 gnd vdd FILL
XFILL_58_DFFSR_182 gnd vdd FILL
XFILL_58_DFFSR_193 gnd vdd FILL
XFILL_32_DFFSR_107 gnd vdd FILL
XFILL_1_DFFSR_120 gnd vdd FILL
XFILL_1_DFFSR_131 gnd vdd FILL
XFILL_21_NOR3X1_3 gnd vdd FILL
XFILL_32_DFFSR_118 gnd vdd FILL
XFILL_32_DFFSR_129 gnd vdd FILL
XFILL_1_DFFSR_142 gnd vdd FILL
XFILL_50_DFFSR_50 gnd vdd FILL
XFILL_1_DFFSR_153 gnd vdd FILL
XFILL_50_DFFSR_61 gnd vdd FILL
XFILL_50_DFFSR_72 gnd vdd FILL
XFILL_1_DFFSR_164 gnd vdd FILL
XFILL_50_DFFSR_83 gnd vdd FILL
XFILL_1_DFFSR_175 gnd vdd FILL
XFILL_21_14 gnd vdd FILL
XFILL_50_DFFSR_94 gnd vdd FILL
XFILL_1_DFFSR_186 gnd vdd FILL
XFILL_1_DFFSR_197 gnd vdd FILL
XFILL_36_DFFSR_106 gnd vdd FILL
XFILL_5_DFFSR_130 gnd vdd FILL
XFILL_36_DFFSR_117 gnd vdd FILL
XFILL_57_1 gnd vdd FILL
XFILL_36_DFFSR_128 gnd vdd FILL
XFILL_5_DFFSR_141 gnd vdd FILL
XFILL_36_DFFSR_139 gnd vdd FILL
XFILL_5_DFFSR_152 gnd vdd FILL
XFILL_5_DFFSR_163 gnd vdd FILL
XFILL_5_DFFSR_174 gnd vdd FILL
XFILL_36_7_0 gnd vdd FILL
XFILL_9_NAND3X1_100 gnd vdd FILL
XFILL_5_DFFSR_185 gnd vdd FILL
XFILL_9_NAND3X1_111 gnd vdd FILL
XFILL_9_NAND3X1_122 gnd vdd FILL
XFILL_5_DFFSR_196 gnd vdd FILL
XFILL_16_MUX2X1_100 gnd vdd FILL
XFILL_9_DFFSR_140 gnd vdd FILL
XFILL_16_MUX2X1_111 gnd vdd FILL
XFILL_4_NOR3X1_4 gnd vdd FILL
XFILL_16_MUX2X1_122 gnd vdd FILL
XFILL_9_DFFSR_151 gnd vdd FILL
XFILL_9_DFFSR_162 gnd vdd FILL
XFILL_13_MUX2X1_60 gnd vdd FILL
XFILL_16_MUX2X1_133 gnd vdd FILL
XFILL_16_MUX2X1_144 gnd vdd FILL
XFILL_13_MUX2X1_71 gnd vdd FILL
XFILL_9_DFFSR_173 gnd vdd FILL
XFILL_30_NOR3X1_1 gnd vdd FILL
XFILL_9_DFFSR_184 gnd vdd FILL
XFILL_13_MUX2X1_82 gnd vdd FILL
XFILL_16_MUX2X1_155 gnd vdd FILL
XFILL_50_2_2 gnd vdd FILL
XFILL_13_MUX2X1_93 gnd vdd FILL
XFILL_1_NOR3X1_20 gnd vdd FILL
XFILL_9_DFFSR_195 gnd vdd FILL
XFILL_1_NOR3X1_31 gnd vdd FILL
XFILL_16_MUX2X1_166 gnd vdd FILL
XFILL_1_NOR3X1_42 gnd vdd FILL
XFILL_16_MUX2X1_177 gnd vdd FILL
XFILL_16_MUX2X1_188 gnd vdd FILL
XFILL_82_DFFSR_207 gnd vdd FILL
XFILL_82_DFFSR_218 gnd vdd FILL
XFILL_82_DFFSR_229 gnd vdd FILL
XFILL_3_DFFSR_5 gnd vdd FILL
XFILL_17_MUX2X1_70 gnd vdd FILL
XFILL_17_MUX2X1_81 gnd vdd FILL
XFILL_17_MUX2X1_92 gnd vdd FILL
XFILL_16_DFFSR_3 gnd vdd FILL
XFILL_5_NOR3X1_30 gnd vdd FILL
XFILL_2_DFFSR_50 gnd vdd FILL
XFILL_5_NOR3X1_41 gnd vdd FILL
XFILL_73_DFFSR_4 gnd vdd FILL
XFILL_5_NOR3X1_52 gnd vdd FILL
XFILL_2_DFFSR_61 gnd vdd FILL
XFILL_86_DFFSR_206 gnd vdd FILL
XFILL_2_DFFSR_72 gnd vdd FILL
XFILL_2_DFFSR_83 gnd vdd FILL
XFILL_86_DFFSR_217 gnd vdd FILL
XFILL_2_DFFSR_94 gnd vdd FILL
XFILL_86_DFFSR_228 gnd vdd FILL
XFILL_21_DFFSR_150 gnd vdd FILL
XFILL_86_DFFSR_239 gnd vdd FILL
XFILL_21_DFFSR_161 gnd vdd FILL
XFILL_21_DFFSR_172 gnd vdd FILL
XFILL_21_DFFSR_183 gnd vdd FILL
XFILL_2_INVX1_101 gnd vdd FILL
XFILL_2_INVX1_112 gnd vdd FILL
XFILL_9_NOR3X1_40 gnd vdd FILL
XFILL_2_INVX1_123 gnd vdd FILL
XFILL_9_NOR3X1_51 gnd vdd FILL
XFILL_21_DFFSR_194 gnd vdd FILL
XFILL_11_BUFX2_9 gnd vdd FILL
XFILL_2_INVX1_134 gnd vdd FILL
XFILL_2_INVX1_145 gnd vdd FILL
XFILL_2_INVX1_156 gnd vdd FILL
XFILL_2_INVX1_167 gnd vdd FILL
XFILL_25_DFFSR_160 gnd vdd FILL
XFILL_2_INVX1_178 gnd vdd FILL
XFILL_25_DFFSR_171 gnd vdd FILL
XFILL_6_INVX1_100 gnd vdd FILL
XFILL_2_INVX1_189 gnd vdd FILL
XFILL_25_DFFSR_182 gnd vdd FILL
XFILL_25_DFFSR_193 gnd vdd FILL
XFILL_6_INVX1_111 gnd vdd FILL
XFILL_6_INVX1_122 gnd vdd FILL
XFILL_23_MUX2X1_190 gnd vdd FILL
XFILL_6_INVX1_133 gnd vdd FILL
XFILL_6_INVX1_144 gnd vdd FILL
XFILL_58_3_2 gnd vdd FILL
XFILL_6_INVX1_155 gnd vdd FILL
XFILL_6_MUX2X1_150 gnd vdd FILL
XFILL_6_MUX2X1_161 gnd vdd FILL
XFILL_6_INVX1_166 gnd vdd FILL
XFILL_38_DFFSR_7 gnd vdd FILL
XFILL_6_INVX1_177 gnd vdd FILL
XFILL_6_INVX1_188 gnd vdd FILL
XFILL_29_DFFSR_170 gnd vdd FILL
XFILL_6_MUX2X1_172 gnd vdd FILL
XFILL_6_MUX2X1_183 gnd vdd FILL
XFILL_29_DFFSR_181 gnd vdd FILL
XFILL_6_INVX1_199 gnd vdd FILL
XFILL_6_MUX2X1_194 gnd vdd FILL
XFILL_29_DFFSR_192 gnd vdd FILL
XFILL_21_NOR3X1_50 gnd vdd FILL
XFILL_2_7_0 gnd vdd FILL
XFILL_27_7_0 gnd vdd FILL
XFILL_0_OAI22X1_7 gnd vdd FILL
XFILL_71_DFFSR_250 gnd vdd FILL
XFILL_71_DFFSR_261 gnd vdd FILL
XFILL_71_DFFSR_272 gnd vdd FILL
XFILL_41_2_2 gnd vdd FILL
XFILL_4_OAI22X1_6 gnd vdd FILL
XFILL_10_BUFX4_3 gnd vdd FILL
XFILL_75_DFFSR_260 gnd vdd FILL
XFILL_30_CLKBUF1_1 gnd vdd FILL
XFILL_75_DFFSR_271 gnd vdd FILL
XFILL_10_6_0 gnd vdd FILL
XFILL_8_OAI22X1_5 gnd vdd FILL
XFILL_79_DFFSR_270 gnd vdd FILL
XFILL_53_DFFSR_206 gnd vdd FILL
XFILL_9_NAND3X1_20 gnd vdd FILL
XFILL_53_DFFSR_217 gnd vdd FILL
XFILL_53_DFFSR_228 gnd vdd FILL
XFILL_9_NAND3X1_31 gnd vdd FILL
XFILL_53_DFFSR_239 gnd vdd FILL
XFILL_9_NAND3X1_42 gnd vdd FILL
XFILL_9_NAND3X1_53 gnd vdd FILL
XFILL_9_NAND3X1_64 gnd vdd FILL
XFILL_15_BUFX4_11 gnd vdd FILL
XFILL_9_NAND3X1_75 gnd vdd FILL
XFILL_15_BUFX4_22 gnd vdd FILL
XFILL_9_NAND3X1_86 gnd vdd FILL
XFILL_80_DFFSR_106 gnd vdd FILL
XFILL_57_DFFSR_205 gnd vdd FILL
XFILL_15_BUFX4_33 gnd vdd FILL
XFILL_9_NAND3X1_97 gnd vdd FILL
XFILL_80_DFFSR_117 gnd vdd FILL
XFILL_15_BUFX4_44 gnd vdd FILL
XFILL_57_DFFSR_216 gnd vdd FILL
XFILL_80_DFFSR_128 gnd vdd FILL
XFILL_15_BUFX4_55 gnd vdd FILL
XFILL_57_DFFSR_227 gnd vdd FILL
XFILL_57_DFFSR_238 gnd vdd FILL
XFILL_80_DFFSR_139 gnd vdd FILL
XFILL_15_BUFX4_66 gnd vdd FILL
XFILL_57_DFFSR_249 gnd vdd FILL
XFILL_15_BUFX4_77 gnd vdd FILL
XFILL_15_BUFX4_88 gnd vdd FILL
XFILL_49_3_2 gnd vdd FILL
XFILL_15_BUFX4_99 gnd vdd FILL
XFILL_84_DFFSR_105 gnd vdd FILL
XFILL_0_DFFSR_209 gnd vdd FILL
XFILL_84_DFFSR_116 gnd vdd FILL
XFILL_84_DFFSR_127 gnd vdd FILL
XFILL_84_DFFSR_138 gnd vdd FILL
XFILL_84_DFFSR_149 gnd vdd FILL
XFILL_2_NAND2X1_11 gnd vdd FILL
XFILL_18_7_0 gnd vdd FILL
XFILL_2_NAND2X1_22 gnd vdd FILL
XFILL_2_NAND2X1_33 gnd vdd FILL
XFILL_2_NAND2X1_44 gnd vdd FILL
XFILL_2_NAND2X1_55 gnd vdd FILL
XFILL_4_DFFSR_208 gnd vdd FILL
XFILL_1_NAND3X1_8 gnd vdd FILL
XFILL_4_DFFSR_219 gnd vdd FILL
XFILL_2_NAND2X1_66 gnd vdd FILL
XFILL_2_NAND2X1_77 gnd vdd FILL
XFILL_0_INVX8_3 gnd vdd FILL
XFILL_2_NAND2X1_88 gnd vdd FILL
XFILL_13_INVX8_1 gnd vdd FILL
XFILL_60_5_0 gnd vdd FILL
XFILL_32_2_2 gnd vdd FILL
XFILL_8_DFFSR_207 gnd vdd FILL
XFILL_10_CLKBUF1_19 gnd vdd FILL
XFILL_5_NAND3X1_7 gnd vdd FILL
XFILL_8_DFFSR_218 gnd vdd FILL
XFILL_8_DFFSR_229 gnd vdd FILL
XFILL_42_DFFSR_260 gnd vdd FILL
XFILL_42_DFFSR_271 gnd vdd FILL
XFILL_9_NAND3X1_6 gnd vdd FILL
XFILL_28_CLKBUF1_10 gnd vdd FILL
XFILL_28_CLKBUF1_21 gnd vdd FILL
XFILL_16_14 gnd vdd FILL
XFILL_28_CLKBUF1_32 gnd vdd FILL
XFILL_55_DFFSR_1 gnd vdd FILL
XFILL_7_BUFX4_10 gnd vdd FILL
XFILL_7_BUFX4_21 gnd vdd FILL
XFILL_7_BUFX4_32 gnd vdd FILL
XFILL_7_BUFX4_43 gnd vdd FILL
XFILL_46_DFFSR_270 gnd vdd FILL
XFILL_7_BUFX4_54 gnd vdd FILL
XFILL_7_BUFX4_65 gnd vdd FILL
XFILL_42_DFFSR_19 gnd vdd FILL
XFILL_7_BUFX4_76 gnd vdd FILL
XFILL_20_DFFSR_206 gnd vdd FILL
XFILL_6_AOI21X1_11 gnd vdd FILL
XFILL_10_NOR2X1_19 gnd vdd FILL
XFILL_20_DFFSR_217 gnd vdd FILL
XFILL_7_BUFX4_87 gnd vdd FILL
XFILL_6_AOI21X1_22 gnd vdd FILL
XFILL_20_DFFSR_228 gnd vdd FILL
XFILL_7_BUFX4_98 gnd vdd FILL
XFILL_6_AOI21X1_33 gnd vdd FILL
XFILL_20_DFFSR_239 gnd vdd FILL
XFILL_6_AOI21X1_44 gnd vdd FILL
XFILL_6_AOI21X1_55 gnd vdd FILL
XFILL_73_DFFSR_170 gnd vdd FILL
XFILL_16_OAI22X1_13 gnd vdd FILL
XFILL_6_AOI21X1_66 gnd vdd FILL
XFILL_16_OAI22X1_24 gnd vdd FILL
XFILL_73_DFFSR_181 gnd vdd FILL
XFILL_16_OAI22X1_35 gnd vdd FILL
XFILL_6_AOI21X1_77 gnd vdd FILL
XFILL_82_DFFSR_18 gnd vdd FILL
XFILL_73_DFFSR_192 gnd vdd FILL
XFILL_24_DFFSR_205 gnd vdd FILL
XFILL_16_OAI22X1_46 gnd vdd FILL
XFILL_82_DFFSR_29 gnd vdd FILL
XFILL_24_DFFSR_216 gnd vdd FILL
XFILL_9_NOR2X1_110 gnd vdd FILL
XFILL_24_DFFSR_227 gnd vdd FILL
XFILL_9_NOR2X1_121 gnd vdd FILL
XFILL_9_NOR2X1_132 gnd vdd FILL
XFILL_24_DFFSR_238 gnd vdd FILL
XFILL_11_DFFSR_18 gnd vdd FILL
XFILL_7_DFFSR_6 gnd vdd FILL
XFILL_9_NOR2X1_143 gnd vdd FILL
XFILL_24_DFFSR_249 gnd vdd FILL
XFILL_11_DFFSR_29 gnd vdd FILL
XFILL_9_NOR2X1_154 gnd vdd FILL
XFILL_0_CLKBUF1_14 gnd vdd FILL
XFILL_0_CLKBUF1_25 gnd vdd FILL
XFILL_77_DFFSR_180 gnd vdd FILL
XFILL_9_NOR2X1_165 gnd vdd FILL
XFILL_77_DFFSR_5 gnd vdd FILL
XFILL_0_CLKBUF1_36 gnd vdd FILL
XFILL_9_NOR2X1_176 gnd vdd FILL
XFILL_77_DFFSR_191 gnd vdd FILL
XFILL_9_NOR2X1_187 gnd vdd FILL
XFILL_51_DFFSR_105 gnd vdd FILL
XFILL_28_DFFSR_204 gnd vdd FILL
XFILL_9_NOR2X1_198 gnd vdd FILL
XFILL_51_DFFSR_116 gnd vdd FILL
XFILL_28_DFFSR_215 gnd vdd FILL
XFILL_51_DFFSR_127 gnd vdd FILL
XFILL_28_DFFSR_226 gnd vdd FILL
XFILL_51_DFFSR_138 gnd vdd FILL
XFILL_28_DFFSR_237 gnd vdd FILL
XFILL_51_DFFSR_17 gnd vdd FILL
XFILL_51_DFFSR_149 gnd vdd FILL
XFILL_28_DFFSR_248 gnd vdd FILL
XFILL_51_DFFSR_28 gnd vdd FILL
XFILL_28_DFFSR_259 gnd vdd FILL
XFILL_51_DFFSR_39 gnd vdd FILL
XFILL_55_DFFSR_104 gnd vdd FILL
XFILL_51_5_0 gnd vdd FILL
XFILL_55_DFFSR_115 gnd vdd FILL
XFILL_55_DFFSR_126 gnd vdd FILL
XFILL_55_DFFSR_137 gnd vdd FILL
XFILL_23_2_2 gnd vdd FILL
XFILL_55_DFFSR_148 gnd vdd FILL
XFILL_55_DFFSR_159 gnd vdd FILL
XFILL_8_MUX2X1_9 gnd vdd FILL
XFILL_20_DFFSR_16 gnd vdd FILL
XFILL_9_MUX2X1_105 gnd vdd FILL
XFILL_59_DFFSR_103 gnd vdd FILL
XFILL_20_DFFSR_27 gnd vdd FILL
XFILL_9_MUX2X1_116 gnd vdd FILL
XFILL_20_DFFSR_38 gnd vdd FILL
XFILL_59_DFFSR_114 gnd vdd FILL
XFILL_11_BUFX4_70 gnd vdd FILL
XFILL_9_MUX2X1_127 gnd vdd FILL
XFILL_59_DFFSR_125 gnd vdd FILL
XFILL_59_DFFSR_136 gnd vdd FILL
XFILL_11_BUFX4_81 gnd vdd FILL
XFILL_9_MUX2X1_138 gnd vdd FILL
XFILL_20_DFFSR_49 gnd vdd FILL
XFILL_9_MUX2X1_149 gnd vdd FILL
XFILL_59_DFFSR_147 gnd vdd FILL
XFILL_11_BUFX4_92 gnd vdd FILL
XFILL_59_DFFSR_158 gnd vdd FILL
XFILL_6_OAI22X1_30 gnd vdd FILL
XFILL_59_DFFSR_169 gnd vdd FILL
XFILL_6_OAI22X1_41 gnd vdd FILL
XFILL_2_DFFSR_107 gnd vdd FILL
XFILL_60_DFFSR_15 gnd vdd FILL
XFILL_60_DFFSR_26 gnd vdd FILL
XFILL_2_DFFSR_118 gnd vdd FILL
XDFFSR_40 DFFSR_40/Q DFFSR_47/CLK DFFSR_79/R vdd DFFSR_40/D gnd vdd DFFSR
XFILL_60_DFFSR_37 gnd vdd FILL
XFILL_2_DFFSR_129 gnd vdd FILL
XFILL_60_DFFSR_48 gnd vdd FILL
XDFFSR_51 INVX1_9/A DFFSR_55/CLK DFFSR_55/R vdd DFFSR_51/D gnd vdd DFFSR
XDFFSR_62 DFFSR_62/Q DFFSR_76/CLK DFFSR_69/R vdd DFFSR_62/D gnd vdd DFFSR
XFILL_60_DFFSR_59 gnd vdd FILL
XDFFSR_73 DFFSR_73/Q DFFSR_73/CLK DFFSR_73/R vdd DFFSR_73/D gnd vdd DFFSR
XDFFSR_84 DFFSR_84/Q DFFSR_84/CLK DFFSR_84/R vdd DFFSR_84/D gnd vdd DFFSR
XDFFSR_95 DFFSR_95/Q DFFSR_99/CLK DFFSR_98/R vdd DFFSR_95/D gnd vdd DFFSR
XFILL_6_DFFSR_106 gnd vdd FILL
XFILL_13_DFFSR_270 gnd vdd FILL
XFILL_6_DFFSR_117 gnd vdd FILL
XFILL_10_MUX2X1_15 gnd vdd FILL
XFILL_3_DFFSR_17 gnd vdd FILL
XFILL_6_DFFSR_128 gnd vdd FILL
XFILL_10_MUX2X1_26 gnd vdd FILL
XFILL_10_MUX2X1_37 gnd vdd FILL
XFILL_3_DFFSR_28 gnd vdd FILL
XFILL_6_DFFSR_139 gnd vdd FILL
XFILL_3_DFFSR_39 gnd vdd FILL
XFILL_1_BUFX4_6 gnd vdd FILL
XFILL_1_AOI21X1_2 gnd vdd FILL
XFILL_10_MUX2X1_48 gnd vdd FILL
XFILL_14_BUFX4_4 gnd vdd FILL
XFILL_10_MUX2X1_59 gnd vdd FILL
XFILL_59_6_0 gnd vdd FILL
XFILL_40_DFFSR_170 gnd vdd FILL
XFILL_6_3_2 gnd vdd FILL
XFILL_5_NAND3X1_130 gnd vdd FILL
XFILL_40_DFFSR_181 gnd vdd FILL
XFILL_5_INVX1_60 gnd vdd FILL
XFILL_14_MUX2X1_14 gnd vdd FILL
XFILL_14_MUX2X1_25 gnd vdd FILL
XFILL_5_INVX1_71 gnd vdd FILL
XFILL_40_DFFSR_192 gnd vdd FILL
XFILL_5_INVX1_82 gnd vdd FILL
XFILL_14_MUX2X1_36 gnd vdd FILL
XFILL_5_INVX1_93 gnd vdd FILL
XFILL_5_AOI21X1_1 gnd vdd FILL
XFILL_14_MUX2X1_47 gnd vdd FILL
XFILL_14_MUX2X1_58 gnd vdd FILL
XFILL_14_MUX2X1_69 gnd vdd FILL
XFILL_12_MUX2X1_3 gnd vdd FILL
XFILL_2_NOR3X1_18 gnd vdd FILL
XFILL_44_DFFSR_180 gnd vdd FILL
XFILL_2_NOR3X1_29 gnd vdd FILL
XFILL_18_MUX2X1_13 gnd vdd FILL
XFILL_44_DFFSR_191 gnd vdd FILL
XFILL_18_MUX2X1_24 gnd vdd FILL
XFILL_18_MUX2X1_35 gnd vdd FILL
XFILL_12_AOI21X1_80 gnd vdd FILL
XFILL_18_MUX2X1_46 gnd vdd FILL
XFILL_18_MUX2X1_57 gnd vdd FILL
XFILL_18_MUX2X1_68 gnd vdd FILL
XFILL_18_MUX2X1_79 gnd vdd FILL
XFILL_6_NOR3X1_17 gnd vdd FILL
XFILL_42_5_0 gnd vdd FILL
XFILL_6_NOR3X1_28 gnd vdd FILL
XFILL_14_2_2 gnd vdd FILL
XFILL_3_BUFX4_80 gnd vdd FILL
XFILL_48_DFFSR_190 gnd vdd FILL
XFILL_6_NOR3X1_39 gnd vdd FILL
XFILL_22_DFFSR_104 gnd vdd FILL
XFILL_3_BUFX4_91 gnd vdd FILL
XFILL_22_DFFSR_115 gnd vdd FILL
XFILL_22_DFFSR_126 gnd vdd FILL
XFILL_22_DFFSR_137 gnd vdd FILL
XFILL_22_DFFSR_148 gnd vdd FILL
XFILL_22_DFFSR_159 gnd vdd FILL
XFILL_26_DFFSR_103 gnd vdd FILL
XFILL_21_MUX2X1_1 gnd vdd FILL
XFILL_26_DFFSR_114 gnd vdd FILL
XFILL_1_NAND3X1_19 gnd vdd FILL
XFILL_26_DFFSR_125 gnd vdd FILL
XFILL_26_DFFSR_136 gnd vdd FILL
XFILL_26_DFFSR_147 gnd vdd FILL
XFILL_26_DFFSR_158 gnd vdd FILL
XINVX1_101 INVX1_101/A gnd NOR3X1_45/A vdd INVX1
XFILL_26_DFFSR_169 gnd vdd FILL
XINVX1_112 INVX1_112/A gnd INVX1_112/Y vdd INVX1
XFILL_5_NOR2X1_4 gnd vdd FILL
XFILL_7_INVX1_109 gnd vdd FILL
XINVX1_123 OAI21X1_9/B gnd INVX1_123/Y vdd INVX1
XINVX1_134 INVX1_134/A gnd INVX1_134/Y vdd INVX1
XINVX1_145 INVX1_145/A gnd NOR3X1_40/A vdd INVX1
XINVX1_156 INVX1_156/A gnd INVX1_156/Y vdd INVX1
XFILL_4_INVX8_4 gnd vdd FILL
XINVX1_167 INVX1_167/A gnd INVX1_167/Y vdd INVX1
XFILL_17_INVX8_2 gnd vdd FILL
XFILL_15_MUX2X1_130 gnd vdd FILL
XINVX1_178 INVX1_178/A gnd INVX1_178/Y vdd INVX1
XINVX1_189 INVX1_189/A gnd INVX1_189/Y vdd INVX1
XFILL_15_MUX2X1_141 gnd vdd FILL
XFILL_29_DFFSR_60 gnd vdd FILL
XFILL_29_DFFSR_71 gnd vdd FILL
XFILL_29_DFFSR_82 gnd vdd FILL
XFILL_22_NOR3X1_15 gnd vdd FILL
XFILL_15_MUX2X1_152 gnd vdd FILL
XFILL_15_MUX2X1_163 gnd vdd FILL
XFILL_29_DFFSR_93 gnd vdd FILL
XFILL_22_NOR3X1_26 gnd vdd FILL
XFILL_15_MUX2X1_174 gnd vdd FILL
XFILL_15_MUX2X1_185 gnd vdd FILL
XFILL_22_NOR3X1_37 gnd vdd FILL
XFILL_22_NOR3X1_48 gnd vdd FILL
XFILL_72_DFFSR_204 gnd vdd FILL
XFILL_4_MUX2X1_2 gnd vdd FILL
XFILL_72_DFFSR_215 gnd vdd FILL
XFILL_72_DFFSR_226 gnd vdd FILL
XFILL_72_DFFSR_237 gnd vdd FILL
XFILL_72_DFFSR_248 gnd vdd FILL
XFILL_69_DFFSR_70 gnd vdd FILL
XFILL_21_DFFSR_4 gnd vdd FILL
XFILL_26_NOR3X1_14 gnd vdd FILL
XFILL_69_DFFSR_81 gnd vdd FILL
XFILL_72_DFFSR_259 gnd vdd FILL
XFILL_69_DFFSR_92 gnd vdd FILL
XFILL_26_NOR3X1_25 gnd vdd FILL
XFILL_26_NOR3X1_36 gnd vdd FILL
XFILL_26_NOR3X1_47 gnd vdd FILL
XFILL_76_DFFSR_203 gnd vdd FILL
XFILL_76_DFFSR_214 gnd vdd FILL
XFILL_59_DFFSR_2 gnd vdd FILL
XFILL_64_1_2 gnd vdd FILL
XFILL_76_DFFSR_225 gnd vdd FILL
XFILL_76_DFFSR_236 gnd vdd FILL
XFILL_1_NOR3X1_8 gnd vdd FILL
XFILL_76_DFFSR_247 gnd vdd FILL
XFILL_0_CLKBUF1_1 gnd vdd FILL
XFILL_76_DFFSR_258 gnd vdd FILL
XFILL_11_DFFSR_180 gnd vdd FILL
XFILL_76_DFFSR_269 gnd vdd FILL
XFILL_11_DFFSR_191 gnd vdd FILL
XFILL_34_3 gnd vdd FILL
XFILL_38_DFFSR_80 gnd vdd FILL
XFILL_33_5_0 gnd vdd FILL
XFILL_38_DFFSR_91 gnd vdd FILL
XFILL_27_2 gnd vdd FILL
XFILL_35_CLKBUF1_9 gnd vdd FILL
XFILL_15_DFFSR_190 gnd vdd FILL
XFILL_78_DFFSR_90 gnd vdd FILL
XFILL_43_DFFSR_8 gnd vdd FILL
XFILL_5_MUX2X1_180 gnd vdd FILL
XFILL_5_MUX2X1_191 gnd vdd FILL
XFILL_1_NOR2X1_109 gnd vdd FILL
XFILL_11_NAND2X1_13 gnd vdd FILL
XFILL_11_NAND2X1_24 gnd vdd FILL
XFILL_11_NAND2X1_35 gnd vdd FILL
XFILL_11_NAND2X1_46 gnd vdd FILL
XFILL_1_OAI21X1_5 gnd vdd FILL
XFILL_11_NAND2X1_57 gnd vdd FILL
XFILL_11_NAND2X1_68 gnd vdd FILL
XFILL_9_OAI22X1_18 gnd vdd FILL
XFILL_11_NAND2X1_79 gnd vdd FILL
XFILL_9_OAI22X1_29 gnd vdd FILL
XFILL_55_1_2 gnd vdd FILL
XFILL_43_DFFSR_203 gnd vdd FILL
XFILL_5_OAI21X1_4 gnd vdd FILL
XFILL_43_DFFSR_214 gnd vdd FILL
XFILL_43_DFFSR_225 gnd vdd FILL
XFILL_2_NOR2X1_40 gnd vdd FILL
XFILL_2_NOR2X1_51 gnd vdd FILL
XFILL_43_DFFSR_236 gnd vdd FILL
XFILL_43_DFFSR_247 gnd vdd FILL
XFILL_8_NAND3X1_50 gnd vdd FILL
XFILL_2_NOR2X1_62 gnd vdd FILL
XFILL_43_DFFSR_258 gnd vdd FILL
XFILL_24_5_0 gnd vdd FILL
XFILL_8_NAND3X1_61 gnd vdd FILL
XFILL_2_NOR2X1_73 gnd vdd FILL
XFILL_43_DFFSR_269 gnd vdd FILL
XFILL_8_NAND3X1_72 gnd vdd FILL
XFILL_2_NOR2X1_84 gnd vdd FILL
XNAND3X1_109 NOR3X1_30/Y NOR2X1_81/Y NOR3X1_28/Y gnd NOR2X1_84/B vdd NAND3X1
XFILL_2_NOR2X1_95 gnd vdd FILL
XFILL_8_NAND3X1_83 gnd vdd FILL
XFILL_47_DFFSR_202 gnd vdd FILL
XFILL_8_NAND3X1_94 gnd vdd FILL
XFILL_70_DFFSR_103 gnd vdd FILL
XFILL_47_DFFSR_213 gnd vdd FILL
XFILL_70_DFFSR_114 gnd vdd FILL
XFILL_5_BUFX4_7 gnd vdd FILL
XFILL_9_OAI21X1_3 gnd vdd FILL
XFILL_70_DFFSR_125 gnd vdd FILL
XFILL_70_DFFSR_136 gnd vdd FILL
XFILL_47_DFFSR_224 gnd vdd FILL
XFILL_47_DFFSR_235 gnd vdd FILL
XFILL_10_OAI22X1_1 gnd vdd FILL
XFILL_6_NOR2X1_50 gnd vdd FILL
XFILL_6_NOR2X1_61 gnd vdd FILL
XFILL_47_DFFSR_246 gnd vdd FILL
XFILL_70_DFFSR_147 gnd vdd FILL
XFILL_70_DFFSR_158 gnd vdd FILL
XFILL_47_DFFSR_257 gnd vdd FILL
XFILL_47_DFFSR_268 gnd vdd FILL
XFILL_70_DFFSR_169 gnd vdd FILL
XFILL_6_NOR2X1_72 gnd vdd FILL
XFILL_6_NOR2X1_83 gnd vdd FILL
XFILL_6_NOR2X1_94 gnd vdd FILL
XFILL_11_AOI22X1_11 gnd vdd FILL
XFILL_74_DFFSR_102 gnd vdd FILL
XFILL_74_DFFSR_113 gnd vdd FILL
XFILL_74_DFFSR_124 gnd vdd FILL
XFILL_74_DFFSR_135 gnd vdd FILL
XFILL_74_DFFSR_146 gnd vdd FILL
XFILL_15_AOI21X1_13 gnd vdd FILL
XFILL_74_DFFSR_157 gnd vdd FILL
XFILL_15_AOI21X1_24 gnd vdd FILL
XFILL_74_DFFSR_168 gnd vdd FILL
XFILL_15_AOI21X1_35 gnd vdd FILL
XFILL_15_AOI21X1_46 gnd vdd FILL
XFILL_74_DFFSR_179 gnd vdd FILL
XFILL_1_NAND2X1_30 gnd vdd FILL
XFILL_78_DFFSR_101 gnd vdd FILL
XFILL_1_NAND2X1_41 gnd vdd FILL
XFILL_1_NAND2X1_52 gnd vdd FILL
XFILL_15_AOI21X1_57 gnd vdd FILL
XFILL_15_AOI21X1_68 gnd vdd FILL
XFILL_1_NAND2X1_63 gnd vdd FILL
XFILL_78_DFFSR_112 gnd vdd FILL
XFILL_12_BUFX4_15 gnd vdd FILL
XFILL_15_AOI21X1_79 gnd vdd FILL
XFILL_78_DFFSR_123 gnd vdd FILL
XFILL_78_DFFSR_134 gnd vdd FILL
XFILL_1_NAND2X1_74 gnd vdd FILL
XFILL_12_BUFX4_26 gnd vdd FILL
XFILL_78_DFFSR_145 gnd vdd FILL
XFILL_12_BUFX4_37 gnd vdd FILL
XFILL_1_NAND2X1_85 gnd vdd FILL
XFILL_78_DFFSR_156 gnd vdd FILL
XFILL_12_BUFX4_48 gnd vdd FILL
XFILL_1_NAND2X1_96 gnd vdd FILL
XFILL_12_BUFX4_59 gnd vdd FILL
XFILL_78_DFFSR_167 gnd vdd FILL
XFILL_78_DFFSR_178 gnd vdd FILL
XFILL_78_DFFSR_189 gnd vdd FILL
XFILL_1_BUFX2_3 gnd vdd FILL
XFILL_7_6_0 gnd vdd FILL
XFILL_6_NAND3X1_120 gnd vdd FILL
XFILL_6_NAND3X1_131 gnd vdd FILL
XFILL_2_NAND2X1_6 gnd vdd FILL
XFILL_60_DFFSR_2 gnd vdd FILL
XFILL_46_1_2 gnd vdd FILL
XFILL_27_CLKBUF1_40 gnd vdd FILL
XFILL_6_INVX1_16 gnd vdd FILL
XFILL_6_NAND2X1_5 gnd vdd FILL
XFILL_10_DFFSR_203 gnd vdd FILL
XFILL_6_INVX1_27 gnd vdd FILL
XFILL_6_INVX1_38 gnd vdd FILL
XFILL_15_5_0 gnd vdd FILL
XFILL_10_DFFSR_214 gnd vdd FILL
XFILL_18_MUX2X1_107 gnd vdd FILL
XFILL_18_MUX2X1_118 gnd vdd FILL
XFILL_7_AND2X2_8 gnd vdd FILL
XFILL_6_INVX1_49 gnd vdd FILL
XFILL_10_DFFSR_225 gnd vdd FILL
XFILL_18_MUX2X1_129 gnd vdd FILL
XFILL_5_AOI21X1_30 gnd vdd FILL
XFILL_10_DFFSR_236 gnd vdd FILL
XFILL_2_MUX2X1_80 gnd vdd FILL
XFILL_5_AOI21X1_41 gnd vdd FILL
XFILL_10_DFFSR_247 gnd vdd FILL
XFILL_2_MUX2X1_91 gnd vdd FILL
XFILL_5_AOI21X1_52 gnd vdd FILL
XFILL_10_DFFSR_258 gnd vdd FILL
XFILL_15_OAI22X1_10 gnd vdd FILL
XFILL_5_AOI21X1_63 gnd vdd FILL
XFILL_10_DFFSR_269 gnd vdd FILL
XFILL_15_OAI22X1_21 gnd vdd FILL
XFILL_5_AOI21X1_74 gnd vdd FILL
XFILL_15_OAI22X1_32 gnd vdd FILL
XFILL_14_DFFSR_202 gnd vdd FILL
XFILL_15_OAI22X1_43 gnd vdd FILL
XFILL_11_NAND3X1_2 gnd vdd FILL
XFILL_14_DFFSR_213 gnd vdd FILL
XFILL_14_DFFSR_224 gnd vdd FILL
XFILL_14_DFFSR_235 gnd vdd FILL
XFILL_8_NOR2X1_140 gnd vdd FILL
XFILL_14_DFFSR_246 gnd vdd FILL
XFILL_25_DFFSR_5 gnd vdd FILL
XDFFSR_107 INVX1_188/A DFFSR_81/CLK DFFSR_82/R vdd DFFSR_107/D gnd vdd DFFSR
XFILL_6_MUX2X1_90 gnd vdd FILL
XFILL_8_NOR2X1_151 gnd vdd FILL
XFILL_14_DFFSR_257 gnd vdd FILL
XFILL_4_BUFX4_14 gnd vdd FILL
XFILL_14_DFFSR_268 gnd vdd FILL
XFILL_8_NOR2X1_162 gnd vdd FILL
XFILL_82_DFFSR_6 gnd vdd FILL
XDFFSR_118 INVX1_180/A CLKBUF1_31/Y DFFSR_2/R vdd DFFSR_118/D gnd vdd DFFSR
XFILL_4_BUFX4_25 gnd vdd FILL
XFILL_8_NOR2X1_173 gnd vdd FILL
XDFFSR_129 INVX1_173/A DFFSR_2/CLK DFFSR_2/R vdd DFFSR_129/D gnd vdd DFFSR
XFILL_18_DFFSR_201 gnd vdd FILL
XFILL_41_DFFSR_102 gnd vdd FILL
XFILL_8_NOR2X1_184 gnd vdd FILL
XFILL_4_BUFX4_36 gnd vdd FILL
XFILL_4_BUFX4_47 gnd vdd FILL
XFILL_18_DFFSR_212 gnd vdd FILL
XFILL_15_NAND3X1_1 gnd vdd FILL
XFILL_8_NOR2X1_195 gnd vdd FILL
XFILL_41_DFFSR_113 gnd vdd FILL
XFILL_41_DFFSR_124 gnd vdd FILL
XFILL_1_INVX2_3 gnd vdd FILL
XFILL_4_BUFX4_58 gnd vdd FILL
XFILL_4_BUFX4_69 gnd vdd FILL
XFILL_41_DFFSR_135 gnd vdd FILL
XFILL_18_DFFSR_223 gnd vdd FILL
XFILL_18_DFFSR_234 gnd vdd FILL
XFILL_41_DFFSR_146 gnd vdd FILL
XFILL_18_DFFSR_245 gnd vdd FILL
XFILL_41_DFFSR_157 gnd vdd FILL
XFILL_18_DFFSR_256 gnd vdd FILL
XFILL_18_DFFSR_267 gnd vdd FILL
XFILL_41_DFFSR_168 gnd vdd FILL
XFILL_41_DFFSR_179 gnd vdd FILL
XFILL_45_DFFSR_101 gnd vdd FILL
XFILL_45_DFFSR_112 gnd vdd FILL
XFILL_45_DFFSR_123 gnd vdd FILL
XFILL_45_DFFSR_134 gnd vdd FILL
XFILL_45_DFFSR_145 gnd vdd FILL
XFILL_45_DFFSR_156 gnd vdd FILL
XFILL_45_DFFSR_167 gnd vdd FILL
XFILL_45_DFFSR_178 gnd vdd FILL
XFILL_8_MUX2X1_102 gnd vdd FILL
XFILL_49_DFFSR_100 gnd vdd FILL
XFILL_45_DFFSR_189 gnd vdd FILL
XFILL_8_MUX2X1_113 gnd vdd FILL
XFILL_49_DFFSR_111 gnd vdd FILL
XFILL_8_MUX2X1_124 gnd vdd FILL
XFILL_49_DFFSR_122 gnd vdd FILL
XFILL_47_DFFSR_9 gnd vdd FILL
XFILL_49_DFFSR_133 gnd vdd FILL
XFILL_8_MUX2X1_135 gnd vdd FILL
XFILL_8_MUX2X1_146 gnd vdd FILL
XFILL_49_DFFSR_144 gnd vdd FILL
XFILL_49_DFFSR_155 gnd vdd FILL
XNOR3X1_18 NOR3X1_18/A NOR3X1_18/B NOR3X1_18/C gnd NOR3X1_18/Y vdd NOR3X1
XFILL_11_AND2X2_2 gnd vdd FILL
XFILL_8_MUX2X1_157 gnd vdd FILL
XFILL_8_MUX2X1_168 gnd vdd FILL
XNOR3X1_29 INVX1_40/Y NOR3X1_29/B NOR3X1_6/C gnd NOR3X1_30/A vdd NOR3X1
XFILL_11_AOI22X1_7 gnd vdd FILL
XFILL_49_DFFSR_166 gnd vdd FILL
XFILL_65_4_0 gnd vdd FILL
XFILL_49_DFFSR_177 gnd vdd FILL
XFILL_8_MUX2X1_179 gnd vdd FILL
XFILL_37_1_2 gnd vdd FILL
XFILL_49_DFFSR_188 gnd vdd FILL
XFILL_49_DFFSR_199 gnd vdd FILL
XFILL_9_OAI21X1_40 gnd vdd FILL
XFILL_15_AOI22X1_6 gnd vdd FILL
XFILL_19_AOI22X1_5 gnd vdd FILL
XFILL_20_0_2 gnd vdd FILL
XFILL_39_DFFSR_14 gnd vdd FILL
XFILL_39_DFFSR_25 gnd vdd FILL
XFILL_39_DFFSR_36 gnd vdd FILL
XFILL_39_DFFSR_47 gnd vdd FILL
XFILL_39_DFFSR_58 gnd vdd FILL
XFILL_39_DFFSR_69 gnd vdd FILL
XFILL_79_DFFSR_13 gnd vdd FILL
XFILL_79_DFFSR_24 gnd vdd FILL
XFILL_79_DFFSR_35 gnd vdd FILL
XFILL_79_DFFSR_46 gnd vdd FILL
XFILL_79_DFFSR_57 gnd vdd FILL
XFILL_79_DFFSR_68 gnd vdd FILL
XFILL_10_NOR2X1_9 gnd vdd FILL
XFILL_79_DFFSR_79 gnd vdd FILL
XFILL_2_INVX1_20 gnd vdd FILL
XFILL_2_INVX1_31 gnd vdd FILL
XFILL_12_DFFSR_101 gnd vdd FILL
XFILL_2_INVX1_42 gnd vdd FILL
XFILL_3_AND2X2_1 gnd vdd FILL
XFILL_2_INVX1_53 gnd vdd FILL
XFILL_12_DFFSR_112 gnd vdd FILL
XFILL_9_BUFX4_8 gnd vdd FILL
XFILL_12_DFFSR_123 gnd vdd FILL
XFILL_12_DFFSR_134 gnd vdd FILL
XFILL_2_INVX1_64 gnd vdd FILL
XFILL_48_DFFSR_12 gnd vdd FILL
XFILL_12_DFFSR_145 gnd vdd FILL
XFILL_2_INVX1_75 gnd vdd FILL
XFILL_2_INVX1_86 gnd vdd FILL
XFILL_48_DFFSR_23 gnd vdd FILL
XFILL_12_DFFSR_156 gnd vdd FILL
XFILL_2_INVX1_97 gnd vdd FILL
XFILL_12_DFFSR_167 gnd vdd FILL
XFILL_48_DFFSR_34 gnd vdd FILL
XFILL_12_DFFSR_178 gnd vdd FILL
XFILL_19_NOR3X1_9 gnd vdd FILL
XFILL_48_DFFSR_45 gnd vdd FILL
XFILL_48_DFFSR_56 gnd vdd FILL
XFILL_16_DFFSR_100 gnd vdd FILL
XFILL_12_DFFSR_189 gnd vdd FILL
XFILL_48_DFFSR_67 gnd vdd FILL
XFILL_48_DFFSR_78 gnd vdd FILL
XFILL_16_DFFSR_111 gnd vdd FILL
XFILL_0_NAND3X1_16 gnd vdd FILL
XFILL_16_DFFSR_122 gnd vdd FILL
XFILL_48_DFFSR_89 gnd vdd FILL
XFILL_56_4_0 gnd vdd FILL
XFILL_16_DFFSR_133 gnd vdd FILL
XFILL_0_NAND3X1_27 gnd vdd FILL
XFILL_16_DFFSR_144 gnd vdd FILL
XFILL_28_1_2 gnd vdd FILL
XFILL_3_1_2 gnd vdd FILL
XFILL_0_NAND3X1_38 gnd vdd FILL
XFILL_16_DFFSR_155 gnd vdd FILL
XFILL_0_NAND3X1_49 gnd vdd FILL
XFILL_16_DFFSR_166 gnd vdd FILL
XFILL_5_CLKBUF1_9 gnd vdd FILL
XFILL_16_DFFSR_177 gnd vdd FILL
XFILL_0_BUFX4_40 gnd vdd FILL
XFILL_4_NAND2X1_18 gnd vdd FILL
XFILL_17_DFFSR_11 gnd vdd FILL
XFILL_16_DFFSR_188 gnd vdd FILL
XFILL_4_NAND2X1_29 gnd vdd FILL
XFILL_0_BUFX4_51 gnd vdd FILL
XFILL_17_DFFSR_22 gnd vdd FILL
XFILL_16_DFFSR_199 gnd vdd FILL
XFILL_17_DFFSR_33 gnd vdd FILL
XFILL_0_BUFX4_62 gnd vdd FILL
XFILL_0_BUFX4_73 gnd vdd FILL
XFILL_0_BUFX4_84 gnd vdd FILL
XFILL_17_DFFSR_44 gnd vdd FILL
XFILL_0_BUFX4_95 gnd vdd FILL
XFILL_17_DFFSR_55 gnd vdd FILL
XFILL_17_DFFSR_66 gnd vdd FILL
XFILL_17_DFFSR_77 gnd vdd FILL
XFILL_1_BUFX4_104 gnd vdd FILL
XFILL_17_DFFSR_88 gnd vdd FILL
XFILL_9_CLKBUF1_8 gnd vdd FILL
XFILL_12_NOR3X1_12 gnd vdd FILL
XFILL_17_DFFSR_99 gnd vdd FILL
XFILL_12_NOR3X1_23 gnd vdd FILL
XFILL_14_MUX2X1_160 gnd vdd FILL
XFILL_57_DFFSR_10 gnd vdd FILL
XFILL_57_DFFSR_21 gnd vdd FILL
XFILL_5_BUFX2_4 gnd vdd FILL
XFILL_14_MUX2X1_171 gnd vdd FILL
XFILL_12_NOR3X1_34 gnd vdd FILL
XFILL_14_MUX2X1_182 gnd vdd FILL
XFILL_57_DFFSR_32 gnd vdd FILL
XFILL_62_DFFSR_201 gnd vdd FILL
XFILL_57_DFFSR_43 gnd vdd FILL
XFILL_28_NOR3X1_7 gnd vdd FILL
XFILL_14_MUX2X1_193 gnd vdd FILL
XFILL_12_NOR3X1_45 gnd vdd FILL
XFILL_62_DFFSR_212 gnd vdd FILL
XFILL_57_DFFSR_54 gnd vdd FILL
XFILL_57_DFFSR_65 gnd vdd FILL
XFILL_62_DFFSR_223 gnd vdd FILL
XFILL_11_0_2 gnd vdd FILL
XFILL_5_BUFX4_103 gnd vdd FILL
XFILL_57_DFFSR_76 gnd vdd FILL
XFILL_62_DFFSR_234 gnd vdd FILL
XFILL_57_DFFSR_87 gnd vdd FILL
XFILL_62_DFFSR_245 gnd vdd FILL
XFILL_16_NOR3X1_11 gnd vdd FILL
XFILL_57_DFFSR_98 gnd vdd FILL
XFILL_62_DFFSR_256 gnd vdd FILL
XFILL_16_NOR3X1_22 gnd vdd FILL
XFILL_62_DFFSR_267 gnd vdd FILL
XFILL_16_NOR3X1_33 gnd vdd FILL
XFILL_66_DFFSR_200 gnd vdd FILL
XFILL_2_NOR2X1_8 gnd vdd FILL
XFILL_16_NOR3X1_44 gnd vdd FILL
XFILL_64_DFFSR_3 gnd vdd FILL
XFILL_66_DFFSR_211 gnd vdd FILL
XFILL_66_DFFSR_222 gnd vdd FILL
XFILL_9_BUFX4_102 gnd vdd FILL
XFILL_26_DFFSR_20 gnd vdd FILL
XFILL_66_DFFSR_233 gnd vdd FILL
XFILL_26_DFFSR_31 gnd vdd FILL
XFILL_26_DFFSR_42 gnd vdd FILL
XFILL_66_DFFSR_244 gnd vdd FILL
XFILL_66_DFFSR_255 gnd vdd FILL
XFILL_26_DFFSR_53 gnd vdd FILL
XFILL_66_DFFSR_266 gnd vdd FILL
XFILL_21_CLKBUF1_7 gnd vdd FILL
XFILL_26_DFFSR_64 gnd vdd FILL
XFILL_26_DFFSR_75 gnd vdd FILL
XFILL_26_DFFSR_86 gnd vdd FILL
XFILL_26_DFFSR_97 gnd vdd FILL
XFILL_8_AOI21X1_18 gnd vdd FILL
XFILL_8_AOI21X1_29 gnd vdd FILL
XFILL_66_DFFSR_30 gnd vdd FILL
XFILL_66_DFFSR_41 gnd vdd FILL
XFILL_1_MUX2X1_6 gnd vdd FILL
XFILL_66_DFFSR_52 gnd vdd FILL
XFILL_66_DFFSR_63 gnd vdd FILL
XFILL_25_CLKBUF1_6 gnd vdd FILL
XFILL_66_DFFSR_74 gnd vdd FILL
XFILL_66_DFFSR_85 gnd vdd FILL
XFILL_66_DFFSR_96 gnd vdd FILL
XFILL_3_NOR2X1_16 gnd vdd FILL
XFILL_3_NOR2X1_27 gnd vdd FILL
XNAND3X1_40 AND2X2_6/A AND2X2_3/B BUFX4_5/Y gnd OAI22X1_32/B vdd NAND3X1
XFILL_3_NOR2X1_38 gnd vdd FILL
XFILL_9_DFFSR_10 gnd vdd FILL
XNAND3X1_51 AND2X2_6/A AND2X2_5/B BUFX4_6/Y gnd INVX1_120/A vdd NAND3X1
XFILL_3_NOR2X1_49 gnd vdd FILL
XNAND3X1_62 BUFX4_57/Y AND2X2_6/B NOR2X1_42/Y gnd OAI22X1_6/B vdd NAND3X1
XFILL_9_DFFSR_21 gnd vdd FILL
XFILL_29_DFFSR_6 gnd vdd FILL
XNAND3X1_73 AND2X2_6/B AND2X2_6/A BUFX4_103/Y gnd OAI22X1_5/B vdd NAND3X1
XFILL_9_DFFSR_32 gnd vdd FILL
XFILL_7_NAND3X1_110 gnd vdd FILL
XFILL_9_DFFSR_43 gnd vdd FILL
XNAND3X1_84 NAND3X1_84/A NOR3X1_13/Y NOR2X1_61/Y gnd NOR3X1_18/C vdd NAND3X1
XFILL_47_4_0 gnd vdd FILL
XFILL_7_NAND3X1_121 gnd vdd FILL
XFILL_9_DFFSR_54 gnd vdd FILL
XFILL_86_DFFSR_7 gnd vdd FILL
XFILL_29_CLKBUF1_5 gnd vdd FILL
XNAND3X1_95 DFFSR_99/Q BUFX4_102/Y NOR2X1_37/Y gnd OAI21X1_16/C vdd NAND3X1
XFILL_7_NAND3X1_132 gnd vdd FILL
XFILL_19_1_2 gnd vdd FILL
XFILL_35_DFFSR_40 gnd vdd FILL
XFILL_9_DFFSR_65 gnd vdd FILL
XFILL_9_DFFSR_76 gnd vdd FILL
XFILL_35_DFFSR_51 gnd vdd FILL
XFILL_7_NOR2X1_15 gnd vdd FILL
XFILL_7_NOR2X1_26 gnd vdd FILL
XFILL_9_DFFSR_87 gnd vdd FILL
XFILL_35_DFFSR_62 gnd vdd FILL
XNOR2X1_40 NOR3X1_49/B NOR2X1_40/B gnd NOR2X1_40/Y vdd NOR2X1
XFILL_5_INVX2_4 gnd vdd FILL
XFILL_9_DFFSR_98 gnd vdd FILL
XNOR2X1_51 INVX1_30/Y NOR2X1_51/B gnd NOR2X1_51/Y vdd NOR2X1
XFILL_7_NOR2X1_37 gnd vdd FILL
XFILL_35_DFFSR_73 gnd vdd FILL
XNOR2X1_62 NOR2X1_62/A NOR2X1_98/B gnd NOR2X1_62/Y vdd NOR2X1
XFILL_7_NOR2X1_48 gnd vdd FILL
XFILL_35_DFFSR_84 gnd vdd FILL
XFILL_7_NOR2X1_59 gnd vdd FILL
XNOR2X1_73 NOR2X1_73/A NOR2X1_73/B gnd NOR2X1_73/Y vdd NOR2X1
XFILL_35_DFFSR_95 gnd vdd FILL
XNOR2X1_84 NOR2X1_84/A NOR2X1_84/B gnd NOR2X1_84/Y vdd NOR2X1
XNOR2X1_95 NOR2X1_95/A NOR2X1_95/B gnd NOR2X1_95/Y vdd NOR2X1
XFILL_0_NOR2X1_106 gnd vdd FILL
XFILL_75_DFFSR_50 gnd vdd FILL
XFILL_0_NOR2X1_117 gnd vdd FILL
XFILL_75_DFFSR_61 gnd vdd FILL
XFILL_0_NOR2X1_128 gnd vdd FILL
XFILL_75_DFFSR_72 gnd vdd FILL
XFILL_75_DFFSR_83 gnd vdd FILL
XFILL_0_NOR2X1_139 gnd vdd FILL
XFILL_15_OAI22X1_9 gnd vdd FILL
XFILL_3_INVX1_2 gnd vdd FILL
XFILL_75_DFFSR_94 gnd vdd FILL
XFILL_11_5 gnd vdd FILL
XFILL_30_3_0 gnd vdd FILL
XFILL_10_NAND2X1_10 gnd vdd FILL
XFILL_10_NAND2X1_21 gnd vdd FILL
XFILL_10_NAND2X1_32 gnd vdd FILL
XFILL_10_NAND2X1_43 gnd vdd FILL
XFILL_15_NOR3X1_2 gnd vdd FILL
XFILL_10_NAND2X1_54 gnd vdd FILL
XFILL_10_NAND2X1_65 gnd vdd FILL
XFILL_19_OAI22X1_8 gnd vdd FILL
XFILL_8_OAI22X1_15 gnd vdd FILL
XFILL_10_NAND2X1_76 gnd vdd FILL
XFILL_10_NAND2X1_87 gnd vdd FILL
XFILL_44_DFFSR_60 gnd vdd FILL
XFILL_8_OAI22X1_26 gnd vdd FILL
XFILL_8_OAI22X1_37 gnd vdd FILL
XFILL_44_DFFSR_71 gnd vdd FILL
XFILL_44_DFFSR_82 gnd vdd FILL
XFILL_8_OAI22X1_48 gnd vdd FILL
XFILL_44_DFFSR_93 gnd vdd FILL
XFILL_33_DFFSR_200 gnd vdd FILL
XFILL_33_DFFSR_211 gnd vdd FILL
XFILL_33_DFFSR_222 gnd vdd FILL
XFILL_33_DFFSR_233 gnd vdd FILL
XFILL_33_DFFSR_244 gnd vdd FILL
XFILL_33_DFFSR_255 gnd vdd FILL
XFILL_84_DFFSR_70 gnd vdd FILL
XFILL_33_DFFSR_266 gnd vdd FILL
XFILL_84_DFFSR_81 gnd vdd FILL
XFILL_84_DFFSR_92 gnd vdd FILL
XFILL_7_NAND3X1_80 gnd vdd FILL
XFILL_7_NAND3X1_91 gnd vdd FILL
XFILL_60_DFFSR_100 gnd vdd FILL
XFILL_37_DFFSR_210 gnd vdd FILL
XFILL_60_DFFSR_111 gnd vdd FILL
XFILL_5_NOR2X1_206 gnd vdd FILL
XFILL_13_DFFSR_70 gnd vdd FILL
XFILL_37_DFFSR_221 gnd vdd FILL
XFILL_60_DFFSR_122 gnd vdd FILL
XFILL_60_DFFSR_133 gnd vdd FILL
XFILL_13_DFFSR_81 gnd vdd FILL
XFILL_13_DFFSR_92 gnd vdd FILL
XFILL_60_DFFSR_144 gnd vdd FILL
XFILL_37_DFFSR_232 gnd vdd FILL
XFILL_37_DFFSR_243 gnd vdd FILL
XFILL_60_DFFSR_155 gnd vdd FILL
XFILL_37_DFFSR_254 gnd vdd FILL
XFILL_60_DFFSR_166 gnd vdd FILL
XFILL_37_DFFSR_265 gnd vdd FILL
XFILL_60_DFFSR_177 gnd vdd FILL
XFILL_3_MUX2X1_12 gnd vdd FILL
XNAND2X1_6 INVX2_1/A NAND2X1_6/B gnd NAND2X1_6/Y vdd NAND2X1
XFILL_3_MUX2X1_23 gnd vdd FILL
XFILL_1_OAI21X1_17 gnd vdd FILL
XFILL_60_DFFSR_188 gnd vdd FILL
XFILL_1_OAI21X1_28 gnd vdd FILL
XFILL_3_MUX2X1_34 gnd vdd FILL
XFILL_3_MUX2X1_45 gnd vdd FILL
XFILL_64_DFFSR_110 gnd vdd FILL
XFILL_60_DFFSR_199 gnd vdd FILL
XFILL_19_CLKBUF1_13 gnd vdd FILL
XFILL_1_OAI21X1_39 gnd vdd FILL
XFILL_19_CLKBUF1_24 gnd vdd FILL
XFILL_64_DFFSR_121 gnd vdd FILL
XFILL_3_MUX2X1_56 gnd vdd FILL
XFILL_53_DFFSR_80 gnd vdd FILL
XFILL_64_DFFSR_132 gnd vdd FILL
XFILL_38_4_0 gnd vdd FILL
XFILL_19_CLKBUF1_35 gnd vdd FILL
XFILL_64_DFFSR_143 gnd vdd FILL
XFILL_53_DFFSR_91 gnd vdd FILL
XFILL_3_MUX2X1_67 gnd vdd FILL
XFILL_64_DFFSR_154 gnd vdd FILL
XFILL_3_MUX2X1_78 gnd vdd FILL
XFILL_14_AOI21X1_10 gnd vdd FILL
XFILL_14_AOI21X1_21 gnd vdd FILL
XFILL_3_MUX2X1_89 gnd vdd FILL
XFILL_14_AOI21X1_32 gnd vdd FILL
XFILL_64_DFFSR_165 gnd vdd FILL
XFILL_7_MUX2X1_11 gnd vdd FILL
XFILL_14_AOI21X1_43 gnd vdd FILL
XFILL_64_DFFSR_176 gnd vdd FILL
XFILL_7_MUX2X1_22 gnd vdd FILL
XFILL_64_DFFSR_187 gnd vdd FILL
XFILL_14_AOI21X1_54 gnd vdd FILL
XFILL_64_DFFSR_198 gnd vdd FILL
XFILL_7_MUX2X1_33 gnd vdd FILL
XFILL_0_NAND2X1_60 gnd vdd FILL
XFILL_7_MUX2X1_44 gnd vdd FILL
XFILL_14_AOI21X1_65 gnd vdd FILL
XFILL_68_DFFSR_120 gnd vdd FILL
XFILL_7_MUX2X1_55 gnd vdd FILL
XFILL_14_AOI21X1_76 gnd vdd FILL
XFILL_0_NAND2X1_71 gnd vdd FILL
XNOR2X1_130 INVX4_1/Y INVX1_174/Y gnd AOI21X1_1/B vdd NOR2X1
XFILL_68_DFFSR_131 gnd vdd FILL
XNOR2X1_141 DFFSR_181/Q AOI21X1_1/B gnd AOI21X1_1/C vdd NOR2X1
XMUX2X1_80 BUFX4_86/Y INVX1_93/Y NOR2X1_28/B gnd MUX2X1_80/Y vdd MUX2X1
XFILL_68_DFFSR_142 gnd vdd FILL
XFILL_7_MUX2X1_66 gnd vdd FILL
XFILL_0_NAND2X1_82 gnd vdd FILL
XNOR2X1_152 INVX2_5/A INVX2_4/Y gnd INVX1_218/A vdd NOR2X1
XFILL_7_MUX2X1_77 gnd vdd FILL
XMUX2X1_91 MUX2X1_91/A BUFX4_96/Y MUX2X1_91/S gnd MUX2X1_91/Y vdd MUX2X1
XFILL_68_DFFSR_153 gnd vdd FILL
XFILL_0_NAND2X1_93 gnd vdd FILL
XFILL_7_MUX2X1_88 gnd vdd FILL
XNOR2X1_163 OAI21X1_46/B INVX1_218/Y gnd INVX1_2/A vdd NOR2X1
XFILL_7_MUX2X1_99 gnd vdd FILL
XNOR2X1_174 INVX4_1/Y INVX1_2/Y gnd MUX2X1_2/S vdd NOR2X1
XFILL_68_DFFSR_164 gnd vdd FILL
XFILL_68_DFFSR_175 gnd vdd FILL
XNOR2X1_185 OAI21X1_46/B INVX1_57/Y gnd INVX1_68/A vdd NOR2X1
XFILL_22_DFFSR_90 gnd vdd FILL
XFILL_68_DFFSR_186 gnd vdd FILL
XNOR2X1_196 INVX4_1/Y INVX1_68/Y gnd NOR2X1_2/B vdd NOR2X1
XFILL_68_DFFSR_197 gnd vdd FILL
XFILL_7_NOR3X1_1 gnd vdd FILL
XFILL_21_3_0 gnd vdd FILL
XMUX2X1_103 NOR3X1_33/A BUFX4_74/Y NAND2X1_16/Y gnd DFFSR_35/D vdd MUX2X1
XMUX2X1_114 BUFX4_68/Y INVX1_156/Y NOR2X1_128/Y gnd DFFSR_144/D vdd MUX2X1
XFILL_5_DFFSR_80 gnd vdd FILL
XFILL_9_CLKBUF1_30 gnd vdd FILL
XMUX2X1_125 BUFX4_99/Y INVX1_169/Y NOR2X1_136/Y gnd DFFSR_133/D vdd MUX2X1
XFILL_5_DFFSR_91 gnd vdd FILL
XMUX2X1_136 BUFX4_66/Y INVX1_180/Y NOR2X1_139/Y gnd DFFSR_118/D vdd MUX2X1
XFILL_23_MUX2X1_20 gnd vdd FILL
XFILL_9_CLKBUF1_41 gnd vdd FILL
XFILL_17_MUX2X1_104 gnd vdd FILL
XFILL_23_MUX2X1_31 gnd vdd FILL
XMUX2X1_147 BUFX4_98/Y INVX1_191/Y NOR2X1_142/Y gnd DFFSR_110/D vdd MUX2X1
XMUX2X1_158 MUX2X1_1/A INVX1_202/Y NOR2X1_156/Y gnd DFFSR_86/D vdd MUX2X1
XFILL_23_MUX2X1_42 gnd vdd FILL
XFILL_23_MUX2X1_53 gnd vdd FILL
XFILL_17_MUX2X1_115 gnd vdd FILL
XFILL_17_MUX2X1_126 gnd vdd FILL
XMUX2X1_169 BUFX4_98/Y INVX1_214/Y NOR2X1_164/Y gnd DFFSR_75/D vdd MUX2X1
XFILL_23_MUX2X1_64 gnd vdd FILL
XFILL_17_MUX2X1_137 gnd vdd FILL
XFILL_23_MUX2X1_75 gnd vdd FILL
XFILL_17_MUX2X1_148 gnd vdd FILL
XFILL_23_MUX2X1_86 gnd vdd FILL
XFILL_4_AOI21X1_60 gnd vdd FILL
XFILL_23_MUX2X1_97 gnd vdd FILL
XFILL_4_AOI21X1_71 gnd vdd FILL
XFILL_9_BUFX2_5 gnd vdd FILL
XFILL_17_MUX2X1_159 gnd vdd FILL
XFILL_14_OAI22X1_40 gnd vdd FILL
XINVX1_10 INVX1_10/A gnd INVX1_10/Y vdd INVX1
XFILL_14_OAI22X1_51 gnd vdd FILL
XINVX1_21 INVX1_21/A gnd NOR3X1_6/A vdd INVX1
XINVX1_32 INVX1_32/A gnd INVX1_32/Y vdd INVX1
XINVX1_43 INVX1_43/A gnd INVX1_43/Y vdd INVX1
XINVX1_54 INVX1_54/A gnd INVX1_54/Y vdd INVX1
XINVX1_65 INVX1_65/A gnd INVX1_65/Y vdd INVX1
XFILL_30_DFFSR_6 gnd vdd FILL
XINVX1_76 INVX1_76/A gnd INVX1_76/Y vdd INVX1
XINVX1_87 INVX1_87/A gnd INVX1_87/Y vdd INVX1
XFILL_29_4_0 gnd vdd FILL
XFILL_4_4_0 gnd vdd FILL
XFILL_7_NOR2X1_170 gnd vdd FILL
XINVX1_98 INVX1_98/A gnd INVX1_98/Y vdd INVX1
XFILL_7_NOR2X1_181 gnd vdd FILL
XFILL_68_DFFSR_4 gnd vdd FILL
XFILL_31_DFFSR_110 gnd vdd FILL
XFILL_7_NOR2X1_192 gnd vdd FILL
XFILL_31_DFFSR_121 gnd vdd FILL
XFILL_31_DFFSR_132 gnd vdd FILL
XFILL_31_DFFSR_143 gnd vdd FILL
XFILL_7_OR2X2_1 gnd vdd FILL
XFILL_31_DFFSR_154 gnd vdd FILL
XFILL_31_DFFSR_165 gnd vdd FILL
XFILL_31_DFFSR_176 gnd vdd FILL
XFILL_31_DFFSR_187 gnd vdd FILL
XFILL_31_DFFSR_198 gnd vdd FILL
XFILL_35_DFFSR_120 gnd vdd FILL
XFILL_35_DFFSR_131 gnd vdd FILL
XFILL_35_DFFSR_142 gnd vdd FILL
XFILL_35_DFFSR_153 gnd vdd FILL
XFILL_35_DFFSR_164 gnd vdd FILL
XFILL_35_DFFSR_175 gnd vdd FILL
XFILL_35_DFFSR_186 gnd vdd FILL
XFILL_12_3_0 gnd vdd FILL
XFILL_35_DFFSR_197 gnd vdd FILL
XFILL_7_MUX2X1_110 gnd vdd FILL
XFILL_7_MUX2X1_121 gnd vdd FILL
XFILL_1_BUFX4_18 gnd vdd FILL
XFILL_1_BUFX4_29 gnd vdd FILL
XFILL_39_DFFSR_130 gnd vdd FILL
XFILL_7_MUX2X1_132 gnd vdd FILL
XFILL_7_MUX2X1_143 gnd vdd FILL
XFILL_39_DFFSR_141 gnd vdd FILL
XFILL_39_DFFSR_152 gnd vdd FILL
XFILL_7_MUX2X1_154 gnd vdd FILL
XFILL_7_MUX2X1_165 gnd vdd FILL
XFILL_39_DFFSR_163 gnd vdd FILL
XFILL_7_MUX2X1_176 gnd vdd FILL
XFILL_39_DFFSR_174 gnd vdd FILL
XFILL_31_NOR3X1_10 gnd vdd FILL
XFILL_7_MUX2X1_187 gnd vdd FILL
XFILL_39_DFFSR_185 gnd vdd FILL
XFILL_31_NOR3X1_21 gnd vdd FILL
XFILL_39_DFFSR_196 gnd vdd FILL
XFILL_31_NOR3X1_32 gnd vdd FILL
XFILL_31_NOR3X1_43 gnd vdd FILL
XFILL_81_DFFSR_210 gnd vdd FILL
XFILL_81_DFFSR_221 gnd vdd FILL
XNOR2X1_9 NOR2X1_9/A NOR2X1_9/B gnd NOR2X1_9/Y vdd NOR2X1
XFILL_81_DFFSR_232 gnd vdd FILL
XFILL_81_DFFSR_243 gnd vdd FILL
XFILL_81_DFFSR_254 gnd vdd FILL
XFILL_81_DFFSR_265 gnd vdd FILL
XFILL_17_DFFSR_109 gnd vdd FILL
XFILL_85_DFFSR_220 gnd vdd FILL
XFILL_12_AOI21X1_5 gnd vdd FILL
XFILL_7_INVX1_3 gnd vdd FILL
XFILL_85_DFFSR_231 gnd vdd FILL
XFILL_85_DFFSR_242 gnd vdd FILL
XFILL_85_DFFSR_253 gnd vdd FILL
XFILL_85_DFFSR_264 gnd vdd FILL
XFILL_85_DFFSR_275 gnd vdd FILL
XFILL_66_6 gnd vdd FILL
XFILL_59_5 gnd vdd FILL
XFILL_1_INVX1_170 gnd vdd FILL
XFILL_8_NAND3X1_100 gnd vdd FILL
XFILL_1_INVX1_181 gnd vdd FILL
XFILL_8_NAND3X1_111 gnd vdd FILL
XFILL_1_INVX1_192 gnd vdd FILL
XFILL_67_DFFSR_19 gnd vdd FILL
XFILL_8_NAND3X1_122 gnd vdd FILL
XFILL_63_7_1 gnd vdd FILL
XFILL_62_2_0 gnd vdd FILL
XFILL_5_INVX1_180 gnd vdd FILL
XFILL_5_INVX1_191 gnd vdd FILL
XFILL_67_DFFSR_209 gnd vdd FILL
XFILL_36_DFFSR_18 gnd vdd FILL
XFILL_36_DFFSR_29 gnd vdd FILL
XAOI21X1_19 BUFX4_76/Y NOR2X1_161/B NOR2X1_160/Y gnd DFFSR_83/D vdd AOI21X1
XFILL_76_DFFSR_17 gnd vdd FILL
XFILL_76_DFFSR_28 gnd vdd FILL
XFILL_76_DFFSR_39 gnd vdd FILL
XFILL_3_NAND2X1_15 gnd vdd FILL
XFILL_19_MUX2X1_7 gnd vdd FILL
XFILL_3_NAND2X1_26 gnd vdd FILL
XFILL_3_NAND2X1_37 gnd vdd FILL
XFILL_3_NAND2X1_48 gnd vdd FILL
XFILL_3_NAND2X1_59 gnd vdd FILL
XFILL_0_AND2X2_5 gnd vdd FILL
XFILL_45_DFFSR_16 gnd vdd FILL
XFILL_45_DFFSR_27 gnd vdd FILL
XFILL_45_DFFSR_38 gnd vdd FILL
XFILL_13_MUX2X1_190 gnd vdd FILL
XFILL_45_DFFSR_49 gnd vdd FILL
XFILL_52_DFFSR_220 gnd vdd FILL
XFILL_52_DFFSR_231 gnd vdd FILL
XFILL_52_DFFSR_242 gnd vdd FILL
XFILL_52_DFFSR_253 gnd vdd FILL
XFILL_85_DFFSR_15 gnd vdd FILL
XFILL_85_DFFSR_26 gnd vdd FILL
XFILL_52_DFFSR_264 gnd vdd FILL
XFILL_12_DFFSR_3 gnd vdd FILL
XFILL_85_DFFSR_37 gnd vdd FILL
XFILL_52_DFFSR_275 gnd vdd FILL
XFILL_85_DFFSR_48 gnd vdd FILL
XFILL_29_CLKBUF1_14 gnd vdd FILL
XFILL_14_DFFSR_15 gnd vdd FILL
XFILL_85_DFFSR_59 gnd vdd FILL
XFILL_29_CLKBUF1_25 gnd vdd FILL
XFILL_14_DFFSR_26 gnd vdd FILL
XFILL_29_CLKBUF1_36 gnd vdd FILL
XFILL_14_DFFSR_37 gnd vdd FILL
XFILL_56_DFFSR_230 gnd vdd FILL
XFILL_54_7_1 gnd vdd FILL
XFILL_56_DFFSR_241 gnd vdd FILL
XFILL_14_DFFSR_48 gnd vdd FILL
XFILL_56_DFFSR_252 gnd vdd FILL
XFILL_14_DFFSR_59 gnd vdd FILL
XFILL_56_DFFSR_263 gnd vdd FILL
XFILL_56_DFFSR_274 gnd vdd FILL
XFILL_53_2_0 gnd vdd FILL
XFILL_11_CLKBUF1_4 gnd vdd FILL
XFILL_54_DFFSR_14 gnd vdd FILL
XFILL_7_AOI21X1_15 gnd vdd FILL
XFILL_54_DFFSR_25 gnd vdd FILL
XFILL_83_DFFSR_130 gnd vdd FILL
XFILL_54_DFFSR_36 gnd vdd FILL
XFILL_7_AOI21X1_26 gnd vdd FILL
XOAI22X1_16 INVX1_47/Y OAI22X1_32/B INVX1_51/Y OAI22X1_32/D gnd NOR2X1_73/A vdd OAI22X1
XOAI22X1_27 MUX2X1_6/A OAI21X1_8/B INVX1_15/Y OAI22X1_36/D gnd NOR2X1_85/B vdd OAI22X1
XFILL_83_DFFSR_141 gnd vdd FILL
XFILL_54_DFFSR_47 gnd vdd FILL
XFILL_83_DFFSR_152 gnd vdd FILL
XFILL_7_AOI21X1_37 gnd vdd FILL
XOAI22X1_38 INVX1_214/Y OAI22X1_48/B INVX1_219/Y OAI22X1_48/D gnd NOR2X1_99/A vdd
+ OAI22X1
XFILL_54_DFFSR_58 gnd vdd FILL
XFILL_7_AOI21X1_48 gnd vdd FILL
XOAI22X1_49 INVX1_197/Y OAI22X1_49/B INVX1_201/Y OAI22X1_49/D gnd NOR2X1_49/A vdd
+ OAI22X1
XFILL_7_AOI21X1_59 gnd vdd FILL
XFILL_54_DFFSR_69 gnd vdd FILL
XFILL_83_DFFSR_163 gnd vdd FILL
XFILL_83_DFFSR_174 gnd vdd FILL
XFILL_15_CLKBUF1_3 gnd vdd FILL
XFILL_17_OAI22X1_17 gnd vdd FILL
XFILL_3_DFFSR_200 gnd vdd FILL
XFILL_17_OAI22X1_28 gnd vdd FILL
XFILL_83_DFFSR_185 gnd vdd FILL
XFILL_3_DFFSR_211 gnd vdd FILL
XFILL_17_OAI22X1_39 gnd vdd FILL
XFILL_83_DFFSR_196 gnd vdd FILL
XFILL_3_DFFSR_222 gnd vdd FILL
XFILL_34_DFFSR_209 gnd vdd FILL
XFILL_3_DFFSR_233 gnd vdd FILL
XFILL_87_DFFSR_140 gnd vdd FILL
XFILL_3_DFFSR_244 gnd vdd FILL
XFILL_87_DFFSR_151 gnd vdd FILL
XFILL_3_DFFSR_255 gnd vdd FILL
XFILL_34_DFFSR_7 gnd vdd FILL
XFILL_23_DFFSR_13 gnd vdd FILL
XFILL_87_DFFSR_162 gnd vdd FILL
XFILL_3_DFFSR_266 gnd vdd FILL
XFILL_1_CLKBUF1_18 gnd vdd FILL
XFILL_23_DFFSR_24 gnd vdd FILL
XFILL_23_DFFSR_35 gnd vdd FILL
XFILL_87_DFFSR_173 gnd vdd FILL
XFILL_19_CLKBUF1_2 gnd vdd FILL
XFILL_87_DFFSR_184 gnd vdd FILL
XFILL_1_CLKBUF1_29 gnd vdd FILL
XFILL_23_DFFSR_46 gnd vdd FILL
XFILL_7_DFFSR_210 gnd vdd FILL
XFILL_23_DFFSR_57 gnd vdd FILL
XFILL_87_DFFSR_195 gnd vdd FILL
XFILL_61_DFFSR_109 gnd vdd FILL
XFILL_38_DFFSR_208 gnd vdd FILL
XFILL_7_DFFSR_221 gnd vdd FILL
XFILL_38_DFFSR_219 gnd vdd FILL
XFILL_23_DFFSR_68 gnd vdd FILL
XFILL_23_DFFSR_79 gnd vdd FILL
XFILL_7_DFFSR_232 gnd vdd FILL
XFILL_7_DFFSR_243 gnd vdd FILL
XFILL_63_DFFSR_12 gnd vdd FILL
XFILL_7_DFFSR_254 gnd vdd FILL
XFILL_7_DFFSR_265 gnd vdd FILL
XFILL_63_DFFSR_23 gnd vdd FILL
XFILL_63_DFFSR_34 gnd vdd FILL
XFILL_63_DFFSR_45 gnd vdd FILL
XFILL_63_DFFSR_56 gnd vdd FILL
XFILL_65_DFFSR_108 gnd vdd FILL
XFILL_63_DFFSR_67 gnd vdd FILL
XFILL_10_OAI21X1_19 gnd vdd FILL
XFILL_65_DFFSR_119 gnd vdd FILL
XFILL_63_DFFSR_78 gnd vdd FILL
XFILL_63_DFFSR_89 gnd vdd FILL
XFILL_8_0_2 gnd vdd FILL
XFILL_6_DFFSR_14 gnd vdd FILL
XFILL_6_DFFSR_25 gnd vdd FILL
XFILL_69_DFFSR_107 gnd vdd FILL
XFILL_32_DFFSR_11 gnd vdd FILL
XFILL_6_DFFSR_36 gnd vdd FILL
XFILL_32_DFFSR_22 gnd vdd FILL
XFILL_6_DFFSR_47 gnd vdd FILL
XFILL_6_DFFSR_58 gnd vdd FILL
XFILL_69_DFFSR_118 gnd vdd FILL
XFILL_69_DFFSR_129 gnd vdd FILL
XFILL_32_DFFSR_33 gnd vdd FILL
XFILL_6_DFFSR_69 gnd vdd FILL
XFILL_0_AOI22X1_5 gnd vdd FILL
XFILL_32_DFFSR_44 gnd vdd FILL
XFILL_32_DFFSR_55 gnd vdd FILL
XFILL_12_OAI21X1_8 gnd vdd FILL
XFILL_7_OAI22X1_12 gnd vdd FILL
XFILL_7_OAI22X1_23 gnd vdd FILL
XFILL_32_DFFSR_66 gnd vdd FILL
XFILL_32_DFFSR_77 gnd vdd FILL
XFILL_7_OAI22X1_34 gnd vdd FILL
XFILL_32_DFFSR_88 gnd vdd FILL
XFILL_7_OAI22X1_45 gnd vdd FILL
XFILL_32_DFFSR_99 gnd vdd FILL
XFILL_0_INVX1_204 gnd vdd FILL
XFILL_72_DFFSR_10 gnd vdd FILL
XFILL_72_DFFSR_21 gnd vdd FILL
XFILL_0_INVX1_215 gnd vdd FILL
XFILL_8_BUFX2_10 gnd vdd FILL
XFILL_45_7_1 gnd vdd FILL
XFILL_72_DFFSR_32 gnd vdd FILL
XFILL_0_INVX1_226 gnd vdd FILL
XFILL_72_DFFSR_43 gnd vdd FILL
XFILL_44_2_0 gnd vdd FILL
XFILL_4_AOI22X1_4 gnd vdd FILL
XFILL_23_DFFSR_230 gnd vdd FILL
XFILL_72_DFFSR_54 gnd vdd FILL
XFILL_23_DFFSR_241 gnd vdd FILL
XFILL_72_DFFSR_65 gnd vdd FILL
XFILL_72_DFFSR_76 gnd vdd FILL
XFILL_23_DFFSR_252 gnd vdd FILL
XFILL_72_DFFSR_87 gnd vdd FILL
XFILL_23_DFFSR_263 gnd vdd FILL
XFILL_23_DFFSR_274 gnd vdd FILL
XFILL_72_DFFSR_98 gnd vdd FILL
XFILL_4_INVX1_203 gnd vdd FILL
XFILL_20_MUX2X1_19 gnd vdd FILL
XFILL_4_INVX1_214 gnd vdd FILL
XFILL_4_INVX1_225 gnd vdd FILL
XFILL_4_NOR2X1_203 gnd vdd FILL
XFILL_50_DFFSR_130 gnd vdd FILL
XFILL_8_AOI22X1_3 gnd vdd FILL
XFILL_50_DFFSR_141 gnd vdd FILL
XFILL_50_DFFSR_152 gnd vdd FILL
XFILL_41_DFFSR_20 gnd vdd FILL
XFILL_27_DFFSR_240 gnd vdd FILL
XFILL_27_DFFSR_251 gnd vdd FILL
XFILL_41_DFFSR_31 gnd vdd FILL
XFILL_12_NOR3X1_6 gnd vdd FILL
XFILL_27_DFFSR_262 gnd vdd FILL
XFILL_41_DFFSR_42 gnd vdd FILL
XFILL_50_DFFSR_163 gnd vdd FILL
XFILL_50_DFFSR_174 gnd vdd FILL
XFILL_27_DFFSR_273 gnd vdd FILL
XFILL_0_OAI21X1_14 gnd vdd FILL
XFILL_41_DFFSR_53 gnd vdd FILL
XFILL_50_DFFSR_185 gnd vdd FILL
XFILL_0_OAI21X1_25 gnd vdd FILL
XFILL_18_CLKBUF1_10 gnd vdd FILL
XFILL_41_DFFSR_64 gnd vdd FILL
XFILL_50_DFFSR_196 gnd vdd FILL
XFILL_0_OAI21X1_36 gnd vdd FILL
XFILL_41_DFFSR_75 gnd vdd FILL
XFILL_18_CLKBUF1_21 gnd vdd FILL
XFILL_41_DFFSR_86 gnd vdd FILL
XFILL_0_OAI21X1_47 gnd vdd FILL
XFILL_18_CLKBUF1_32 gnd vdd FILL
XFILL_41_DFFSR_97 gnd vdd FILL
XFILL_54_DFFSR_140 gnd vdd FILL
XFILL_54_DFFSR_151 gnd vdd FILL
XFILL_54_DFFSR_162 gnd vdd FILL
XFILL_81_DFFSR_30 gnd vdd FILL
XFILL_81_DFFSR_41 gnd vdd FILL
XFILL_13_AOI21X1_40 gnd vdd FILL
XFILL_54_DFFSR_173 gnd vdd FILL
XFILL_81_DFFSR_52 gnd vdd FILL
XFILL_54_DFFSR_184 gnd vdd FILL
XFILL_13_AOI21X1_51 gnd vdd FILL
XFILL_81_DFFSR_63 gnd vdd FILL
XFILL_54_DFFSR_195 gnd vdd FILL
XFILL_13_AOI21X1_62 gnd vdd FILL
XFILL_81_DFFSR_74 gnd vdd FILL
XFILL_10_DFFSR_30 gnd vdd FILL
XFILL_13_AOI21X1_73 gnd vdd FILL
XFILL_81_DFFSR_85 gnd vdd FILL
XFILL_10_DFFSR_41 gnd vdd FILL
XFILL_81_DFFSR_96 gnd vdd FILL
XFILL_10_DFFSR_52 gnd vdd FILL
XFILL_10_DFFSR_63 gnd vdd FILL
XFILL_58_DFFSR_150 gnd vdd FILL
XFILL_8_NOR2X1_1 gnd vdd FILL
XFILL_58_DFFSR_161 gnd vdd FILL
XFILL_10_DFFSR_74 gnd vdd FILL
XFILL_10_DFFSR_85 gnd vdd FILL
XFILL_58_DFFSR_172 gnd vdd FILL
XFILL_10_DFFSR_96 gnd vdd FILL
XFILL_58_DFFSR_183 gnd vdd FILL
XFILL_58_DFFSR_194 gnd vdd FILL
XFILL_1_DFFSR_110 gnd vdd FILL
XFILL_32_DFFSR_108 gnd vdd FILL
XFILL_1_DFFSR_121 gnd vdd FILL
XFILL_50_DFFSR_40 gnd vdd FILL
XFILL_1_DFFSR_132 gnd vdd FILL
XFILL_8_1 gnd vdd FILL
XFILL_32_DFFSR_119 gnd vdd FILL
XFILL_21_NOR3X1_4 gnd vdd FILL
XFILL_50_DFFSR_51 gnd vdd FILL
XFILL_1_DFFSR_143 gnd vdd FILL
XFILL_1_DFFSR_154 gnd vdd FILL
XFILL_50_DFFSR_62 gnd vdd FILL
XFILL_1_DFFSR_165 gnd vdd FILL
XFILL_50_DFFSR_73 gnd vdd FILL
XFILL_21_15 gnd vdd FILL
XFILL_50_DFFSR_84 gnd vdd FILL
XFILL_1_DFFSR_176 gnd vdd FILL
XFILL_50_DFFSR_95 gnd vdd FILL
XFILL_1_DFFSR_187 gnd vdd FILL
XFILL_1_DFFSR_198 gnd vdd FILL
XFILL_36_DFFSR_107 gnd vdd FILL
XFILL_5_DFFSR_120 gnd vdd FILL
XFILL_5_DFFSR_131 gnd vdd FILL
XFILL_36_DFFSR_118 gnd vdd FILL
XFILL_57_2 gnd vdd FILL
XFILL_5_DFFSR_142 gnd vdd FILL
XFILL_36_DFFSR_129 gnd vdd FILL
XFILL_5_DFFSR_153 gnd vdd FILL
XFILL_51_DFFSR_1 gnd vdd FILL
XFILL_5_DFFSR_164 gnd vdd FILL
XFILL_5_DFFSR_175 gnd vdd FILL
XFILL_9_NAND3X1_101 gnd vdd FILL
XFILL_36_7_1 gnd vdd FILL
XFILL_5_DFFSR_186 gnd vdd FILL
XFILL_9_NAND3X1_112 gnd vdd FILL
XFILL_5_DFFSR_197 gnd vdd FILL
XFILL_9_NAND3X1_123 gnd vdd FILL
XFILL_35_2_0 gnd vdd FILL
XFILL_9_DFFSR_130 gnd vdd FILL
XFILL_16_MUX2X1_101 gnd vdd FILL
XFILL_16_MUX2X1_112 gnd vdd FILL
XFILL_9_DFFSR_141 gnd vdd FILL
XFILL_9_DFFSR_152 gnd vdd FILL
XFILL_13_MUX2X1_50 gnd vdd FILL
XFILL_4_NOR3X1_5 gnd vdd FILL
XFILL_16_MUX2X1_123 gnd vdd FILL
XFILL_9_DFFSR_163 gnd vdd FILL
XFILL_13_MUX2X1_61 gnd vdd FILL
XFILL_30_NOR3X1_2 gnd vdd FILL
XFILL_16_MUX2X1_134 gnd vdd FILL
XFILL_9_DFFSR_174 gnd vdd FILL
XFILL_16_MUX2X1_145 gnd vdd FILL
XFILL_1_NOR3X1_10 gnd vdd FILL
XFILL_13_MUX2X1_72 gnd vdd FILL
XFILL_16_MUX2X1_156 gnd vdd FILL
XFILL_13_MUX2X1_83 gnd vdd FILL
XFILL_9_DFFSR_185 gnd vdd FILL
XFILL_1_NOR3X1_21 gnd vdd FILL
XFILL_13_MUX2X1_94 gnd vdd FILL
XFILL_1_NOR3X1_32 gnd vdd FILL
XFILL_9_DFFSR_196 gnd vdd FILL
XFILL_16_MUX2X1_167 gnd vdd FILL
XFILL_16_MUX2X1_178 gnd vdd FILL
XFILL_1_NOR3X1_43 gnd vdd FILL
XFILL_16_MUX2X1_189 gnd vdd FILL
XFILL_82_DFFSR_208 gnd vdd FILL
XFILL_82_DFFSR_219 gnd vdd FILL
XFILL_17_MUX2X1_60 gnd vdd FILL
XFILL_17_MUX2X1_71 gnd vdd FILL
XFILL_3_DFFSR_6 gnd vdd FILL
XFILL_17_MUX2X1_82 gnd vdd FILL
XFILL_5_NOR3X1_20 gnd vdd FILL
XFILL_16_DFFSR_4 gnd vdd FILL
XFILL_2_DFFSR_40 gnd vdd FILL
XFILL_17_MUX2X1_93 gnd vdd FILL
XFILL_5_NOR3X1_31 gnd vdd FILL
XFILL_2_DFFSR_51 gnd vdd FILL
XFILL_5_NOR3X1_42 gnd vdd FILL
XFILL_73_DFFSR_5 gnd vdd FILL
XFILL_2_DFFSR_62 gnd vdd FILL
XFILL_2_DFFSR_73 gnd vdd FILL
XFILL_86_DFFSR_207 gnd vdd FILL
XFILL_2_DFFSR_84 gnd vdd FILL
XFILL_86_DFFSR_218 gnd vdd FILL
XFILL_2_DFFSR_95 gnd vdd FILL
XFILL_21_DFFSR_140 gnd vdd FILL
XFILL_86_DFFSR_229 gnd vdd FILL
XFILL_21_DFFSR_151 gnd vdd FILL
XFILL_21_DFFSR_162 gnd vdd FILL
XFILL_2_INVX1_102 gnd vdd FILL
XFILL_21_DFFSR_173 gnd vdd FILL
XFILL_9_NOR3X1_30 gnd vdd FILL
XFILL_21_DFFSR_184 gnd vdd FILL
XFILL_9_NOR3X1_41 gnd vdd FILL
XFILL_2_INVX1_113 gnd vdd FILL
XFILL_21_DFFSR_195 gnd vdd FILL
XFILL_9_NOR3X1_52 gnd vdd FILL
XFILL_2_INVX1_124 gnd vdd FILL
XFILL_2_INVX1_135 gnd vdd FILL
XFILL_2_INVX1_146 gnd vdd FILL
XFILL_2_INVX1_157 gnd vdd FILL
XFILL_25_DFFSR_150 gnd vdd FILL
XFILL_25_DFFSR_161 gnd vdd FILL
XFILL_2_INVX1_168 gnd vdd FILL
XFILL_2_INVX1_179 gnd vdd FILL
XFILL_25_DFFSR_172 gnd vdd FILL
XFILL_6_INVX1_101 gnd vdd FILL
XFILL_6_INVX1_112 gnd vdd FILL
XFILL_25_DFFSR_183 gnd vdd FILL
XFILL_4_NAND3X1_130 gnd vdd FILL
XFILL_25_DFFSR_194 gnd vdd FILL
XFILL_6_INVX1_123 gnd vdd FILL
XFILL_23_MUX2X1_180 gnd vdd FILL
XFILL_6_INVX1_134 gnd vdd FILL
XFILL_23_MUX2X1_191 gnd vdd FILL
XFILL_6_INVX1_145 gnd vdd FILL
XFILL_6_MUX2X1_140 gnd vdd FILL
XFILL_6_INVX1_156 gnd vdd FILL
XFILL_38_DFFSR_8 gnd vdd FILL
XFILL_6_MUX2X1_151 gnd vdd FILL
XFILL_29_DFFSR_160 gnd vdd FILL
XFILL_6_INVX1_167 gnd vdd FILL
XFILL_6_MUX2X1_162 gnd vdd FILL
XFILL_6_MUX2X1_173 gnd vdd FILL
XFILL_29_DFFSR_171 gnd vdd FILL
XFILL_6_INVX1_178 gnd vdd FILL
XFILL_6_INVX1_189 gnd vdd FILL
XFILL_6_MUX2X1_184 gnd vdd FILL
XFILL_29_DFFSR_182 gnd vdd FILL
XFILL_29_DFFSR_193 gnd vdd FILL
XFILL_21_NOR3X1_40 gnd vdd FILL
XFILL_27_7_1 gnd vdd FILL
XFILL_21_NOR3X1_51 gnd vdd FILL
XFILL_2_7_1 gnd vdd FILL
XFILL_0_OAI22X1_8 gnd vdd FILL
XFILL_26_2_0 gnd vdd FILL
XFILL_1_2_0 gnd vdd FILL
XFILL_71_DFFSR_240 gnd vdd FILL
XFILL_71_DFFSR_251 gnd vdd FILL
XFILL_71_DFFSR_262 gnd vdd FILL
XFILL_71_DFFSR_273 gnd vdd FILL
XFILL_25_NOR3X1_50 gnd vdd FILL
XFILL_4_OAI22X1_7 gnd vdd FILL
XFILL_10_BUFX4_4 gnd vdd FILL
XFILL_75_DFFSR_250 gnd vdd FILL
XFILL_75_DFFSR_261 gnd vdd FILL
XFILL_75_DFFSR_272 gnd vdd FILL
XFILL_30_CLKBUF1_2 gnd vdd FILL
XFILL_10_6_1 gnd vdd FILL
XFILL_8_OAI22X1_6 gnd vdd FILL
XFILL_79_DFFSR_260 gnd vdd FILL
XFILL_79_DFFSR_271 gnd vdd FILL
XFILL_34_CLKBUF1_1 gnd vdd FILL
XFILL_53_DFFSR_207 gnd vdd FILL
XFILL_53_DFFSR_218 gnd vdd FILL
XFILL_9_NAND3X1_10 gnd vdd FILL
XFILL_9_NAND3X1_21 gnd vdd FILL
XFILL_9_NAND3X1_32 gnd vdd FILL
XFILL_53_DFFSR_229 gnd vdd FILL
XFILL_9_NAND3X1_43 gnd vdd FILL
XFILL_9_NAND3X1_54 gnd vdd FILL
XFILL_15_BUFX4_12 gnd vdd FILL
XFILL_9_NAND3X1_65 gnd vdd FILL
XFILL_9_NAND3X1_76 gnd vdd FILL
XFILL_15_BUFX4_23 gnd vdd FILL
XFILL_9_NAND3X1_87 gnd vdd FILL
XFILL_9_3_0 gnd vdd FILL
XFILL_57_DFFSR_206 gnd vdd FILL
XFILL_80_DFFSR_107 gnd vdd FILL
XFILL_15_BUFX4_34 gnd vdd FILL
XFILL_9_NAND3X1_98 gnd vdd FILL
XFILL_15_BUFX4_45 gnd vdd FILL
XFILL_57_DFFSR_217 gnd vdd FILL
XFILL_80_DFFSR_118 gnd vdd FILL
XFILL_57_DFFSR_228 gnd vdd FILL
XFILL_80_DFFSR_129 gnd vdd FILL
XFILL_15_BUFX4_56 gnd vdd FILL
XFILL_15_BUFX4_67 gnd vdd FILL
XFILL_15_BUFX4_78 gnd vdd FILL
XFILL_57_DFFSR_239 gnd vdd FILL
XFILL_15_BUFX4_89 gnd vdd FILL
XFILL_84_DFFSR_106 gnd vdd FILL
XFILL_84_DFFSR_117 gnd vdd FILL
XFILL_84_DFFSR_128 gnd vdd FILL
XFILL_84_DFFSR_139 gnd vdd FILL
XFILL_18_7_1 gnd vdd FILL
XFILL_2_NAND2X1_12 gnd vdd FILL
XFILL_2_NAND2X1_23 gnd vdd FILL
XFILL_17_2_0 gnd vdd FILL
XFILL_2_NAND2X1_34 gnd vdd FILL
XFILL_4_DFFSR_209 gnd vdd FILL
XFILL_2_NAND2X1_45 gnd vdd FILL
XFILL_1_NAND3X1_9 gnd vdd FILL
XFILL_2_NAND2X1_56 gnd vdd FILL
XFILL_2_NAND2X1_67 gnd vdd FILL
XFILL_2_NAND2X1_78 gnd vdd FILL
XFILL_0_INVX8_4 gnd vdd FILL
XFILL_2_NAND2X1_89 gnd vdd FILL
XFILL_13_INVX8_2 gnd vdd FILL
XFILL_60_5_1 gnd vdd FILL
XFILL_8_DFFSR_208 gnd vdd FILL
XFILL_8_DFFSR_219 gnd vdd FILL
XFILL_5_NAND3X1_8 gnd vdd FILL
XFILL_42_DFFSR_250 gnd vdd FILL
XFILL_42_DFFSR_261 gnd vdd FILL
XFILL_42_DFFSR_272 gnd vdd FILL
XFILL_9_NAND3X1_7 gnd vdd FILL
XFILL_28_CLKBUF1_11 gnd vdd FILL
XFILL_28_CLKBUF1_22 gnd vdd FILL
XFILL_16_15 gnd vdd FILL
XFILL_28_CLKBUF1_33 gnd vdd FILL
XFILL_55_DFFSR_2 gnd vdd FILL
XFILL_7_BUFX4_11 gnd vdd FILL
XFILL_7_BUFX4_22 gnd vdd FILL
XFILL_7_BUFX4_33 gnd vdd FILL
XFILL_2_AOI22X1_10 gnd vdd FILL
XFILL_7_BUFX4_44 gnd vdd FILL
XFILL_46_DFFSR_260 gnd vdd FILL
XFILL_46_DFFSR_271 gnd vdd FILL
XFILL_7_BUFX4_55 gnd vdd FILL
XFILL_7_BUFX4_66 gnd vdd FILL
XFILL_20_DFFSR_207 gnd vdd FILL
XFILL_7_BUFX4_77 gnd vdd FILL
XFILL_6_AOI21X1_12 gnd vdd FILL
XFILL_20_DFFSR_218 gnd vdd FILL
XFILL_7_BUFX4_88 gnd vdd FILL
XFILL_7_BUFX4_99 gnd vdd FILL
XFILL_6_AOI21X1_23 gnd vdd FILL
XFILL_20_DFFSR_229 gnd vdd FILL
XFILL_6_AOI21X1_34 gnd vdd FILL
XFILL_73_DFFSR_160 gnd vdd FILL
XFILL_6_AOI21X1_45 gnd vdd FILL
XFILL_16_OAI22X1_14 gnd vdd FILL
XFILL_6_AOI21X1_56 gnd vdd FILL
XFILL_6_AOI21X1_67 gnd vdd FILL
XFILL_73_DFFSR_171 gnd vdd FILL
XFILL_6_AOI21X1_78 gnd vdd FILL
XFILL_16_OAI22X1_25 gnd vdd FILL
XFILL_73_DFFSR_182 gnd vdd FILL
XFILL_82_DFFSR_19 gnd vdd FILL
XFILL_73_DFFSR_193 gnd vdd FILL
XFILL_16_OAI22X1_36 gnd vdd FILL
XFILL_24_DFFSR_206 gnd vdd FILL
XFILL_16_OAI22X1_47 gnd vdd FILL
XFILL_9_NOR2X1_100 gnd vdd FILL
XFILL_24_DFFSR_217 gnd vdd FILL
XFILL_9_NOR2X1_111 gnd vdd FILL
XFILL_24_DFFSR_228 gnd vdd FILL
XFILL_9_NOR2X1_122 gnd vdd FILL
XFILL_11_DFFSR_19 gnd vdd FILL
XFILL_9_NOR2X1_133 gnd vdd FILL
XFILL_24_DFFSR_239 gnd vdd FILL
XFILL_7_DFFSR_7 gnd vdd FILL
XFILL_9_NOR2X1_144 gnd vdd FILL
XFILL_77_DFFSR_170 gnd vdd FILL
XFILL_9_NOR2X1_155 gnd vdd FILL
XFILL_0_CLKBUF1_15 gnd vdd FILL
XFILL_9_NOR2X1_166 gnd vdd FILL
XFILL_0_CLKBUF1_26 gnd vdd FILL
XFILL_77_DFFSR_181 gnd vdd FILL
XFILL_77_DFFSR_6 gnd vdd FILL
XFILL_9_NOR2X1_177 gnd vdd FILL
XFILL_77_DFFSR_192 gnd vdd FILL
XFILL_0_CLKBUF1_37 gnd vdd FILL
XFILL_51_DFFSR_106 gnd vdd FILL
XFILL_28_DFFSR_205 gnd vdd FILL
XFILL_9_NOR2X1_188 gnd vdd FILL
XFILL_9_NOR2X1_199 gnd vdd FILL
XFILL_28_DFFSR_216 gnd vdd FILL
XFILL_51_DFFSR_117 gnd vdd FILL
XFILL_28_DFFSR_227 gnd vdd FILL
XFILL_51_DFFSR_128 gnd vdd FILL
XFILL_15_NAND3X1_90 gnd vdd FILL
XFILL_51_DFFSR_139 gnd vdd FILL
XFILL_28_DFFSR_238 gnd vdd FILL
XFILL_51_DFFSR_18 gnd vdd FILL
XFILL_28_DFFSR_249 gnd vdd FILL
XFILL_51_DFFSR_29 gnd vdd FILL
XFILL_55_DFFSR_105 gnd vdd FILL
XFILL_51_5_1 gnd vdd FILL
XFILL_55_DFFSR_116 gnd vdd FILL
XFILL_55_DFFSR_127 gnd vdd FILL
XFILL_55_DFFSR_138 gnd vdd FILL
XFILL_55_DFFSR_149 gnd vdd FILL
XFILL_50_0_0 gnd vdd FILL
XFILL_59_DFFSR_104 gnd vdd FILL
XFILL_9_MUX2X1_106 gnd vdd FILL
XFILL_20_DFFSR_17 gnd vdd FILL
XFILL_9_MUX2X1_117 gnd vdd FILL
XFILL_20_DFFSR_28 gnd vdd FILL
XFILL_59_DFFSR_115 gnd vdd FILL
XFILL_11_BUFX4_60 gnd vdd FILL
XFILL_20_DFFSR_39 gnd vdd FILL
XFILL_9_MUX2X1_128 gnd vdd FILL
XFILL_11_BUFX4_71 gnd vdd FILL
XFILL_59_DFFSR_126 gnd vdd FILL
XFILL_59_DFFSR_137 gnd vdd FILL
XFILL_9_MUX2X1_139 gnd vdd FILL
XFILL_11_BUFX4_82 gnd vdd FILL
XFILL_59_DFFSR_148 gnd vdd FILL
XFILL_11_BUFX4_93 gnd vdd FILL
XFILL_6_OAI22X1_20 gnd vdd FILL
XFILL_59_DFFSR_159 gnd vdd FILL
XFILL_6_OAI22X1_31 gnd vdd FILL
XFILL_6_OAI22X1_42 gnd vdd FILL
XFILL_60_DFFSR_16 gnd vdd FILL
XFILL_2_DFFSR_108 gnd vdd FILL
XDFFSR_30 DFFSR_30/Q DFFSR_88/CLK DFFSR_4/R vdd DFFSR_30/D gnd vdd DFFSR
XFILL_60_DFFSR_27 gnd vdd FILL
XFILL_2_DFFSR_119 gnd vdd FILL
XFILL_60_DFFSR_38 gnd vdd FILL
XDFFSR_41 INVX1_17/A DFFSR_56/CLK DFFSR_42/R vdd MUX2X1_4/Y gnd vdd DFFSR
XFILL_60_DFFSR_49 gnd vdd FILL
XDFFSR_52 INVX1_10/A DFFSR_52/CLK DFFSR_56/R vdd DFFSR_52/D gnd vdd DFFSR
XDFFSR_63 DFFSR_63/Q DFFSR_97/CLK DFFSR_69/R vdd DFFSR_63/D gnd vdd DFFSR
XDFFSR_74 DFFSR_74/Q DFFSR_76/CLK DFFSR_97/R vdd DFFSR_74/D gnd vdd DFFSR
XDFFSR_85 DFFSR_85/Q DFFSR_93/CLK DFFSR_89/R vdd DFFSR_85/D gnd vdd DFFSR
XDFFSR_96 DFFSR_96/Q CLKBUF1_8/Y DFFSR_96/R vdd DFFSR_96/D gnd vdd DFFSR
XFILL_13_DFFSR_260 gnd vdd FILL
XFILL_6_DFFSR_107 gnd vdd FILL
XFILL_13_DFFSR_271 gnd vdd FILL
XFILL_10_MUX2X1_16 gnd vdd FILL
XFILL_6_DFFSR_118 gnd vdd FILL
XFILL_6_DFFSR_129 gnd vdd FILL
XFILL_3_DFFSR_18 gnd vdd FILL
XFILL_10_MUX2X1_27 gnd vdd FILL
XFILL_3_NOR2X1_200 gnd vdd FILL
XFILL_3_DFFSR_29 gnd vdd FILL
XFILL_10_MUX2X1_38 gnd vdd FILL
XFILL_1_AOI21X1_3 gnd vdd FILL
XFILL_10_MUX2X1_49 gnd vdd FILL
XFILL_1_BUFX4_7 gnd vdd FILL
XFILL_14_BUFX4_5 gnd vdd FILL
XFILL_40_DFFSR_160 gnd vdd FILL
XFILL_59_6_1 gnd vdd FILL
XFILL_5_NAND3X1_120 gnd vdd FILL
XFILL_17_DFFSR_270 gnd vdd FILL
XFILL_5_INVX1_50 gnd vdd FILL
XFILL_40_DFFSR_171 gnd vdd FILL
XFILL_5_NAND3X1_131 gnd vdd FILL
XFILL_5_INVX1_61 gnd vdd FILL
XFILL_14_MUX2X1_15 gnd vdd FILL
XFILL_40_DFFSR_182 gnd vdd FILL
XFILL_58_1_0 gnd vdd FILL
XFILL_5_INVX1_72 gnd vdd FILL
XFILL_40_DFFSR_193 gnd vdd FILL
XFILL_14_MUX2X1_26 gnd vdd FILL
XFILL_5_INVX1_83 gnd vdd FILL
XFILL_14_MUX2X1_37 gnd vdd FILL
XFILL_5_INVX1_94 gnd vdd FILL
XFILL_5_AOI21X1_2 gnd vdd FILL
XFILL_14_MUX2X1_48 gnd vdd FILL
XFILL_14_MUX2X1_59 gnd vdd FILL
XFILL_17_CLKBUF1_40 gnd vdd FILL
XFILL_12_MUX2X1_4 gnd vdd FILL
XFILL_2_NOR3X1_19 gnd vdd FILL
XFILL_44_DFFSR_170 gnd vdd FILL
XFILL_18_MUX2X1_14 gnd vdd FILL
XFILL_44_DFFSR_181 gnd vdd FILL
XFILL_44_DFFSR_192 gnd vdd FILL
XFILL_18_MUX2X1_25 gnd vdd FILL
XFILL_12_AOI21X1_70 gnd vdd FILL
XFILL_18_MUX2X1_36 gnd vdd FILL
XFILL_12_AOI21X1_81 gnd vdd FILL
XFILL_18_MUX2X1_47 gnd vdd FILL
XFILL_9_AOI21X1_1 gnd vdd FILL
XFILL_18_MUX2X1_58 gnd vdd FILL
XFILL_18_MUX2X1_69 gnd vdd FILL
XFILL_42_5_1 gnd vdd FILL
XFILL_6_NOR3X1_18 gnd vdd FILL
XFILL_6_NOR3X1_29 gnd vdd FILL
XFILL_48_DFFSR_180 gnd vdd FILL
XFILL_3_BUFX4_70 gnd vdd FILL
XFILL_3_BUFX4_81 gnd vdd FILL
XFILL_22_DFFSR_105 gnd vdd FILL
XFILL_41_0_0 gnd vdd FILL
XFILL_48_DFFSR_191 gnd vdd FILL
XFILL_3_BUFX4_92 gnd vdd FILL
XFILL_22_DFFSR_116 gnd vdd FILL
XFILL_10_BUFX2_1 gnd vdd FILL
XFILL_22_DFFSR_127 gnd vdd FILL
XFILL_22_DFFSR_138 gnd vdd FILL
XFILL_22_DFFSR_149 gnd vdd FILL
XFILL_26_DFFSR_104 gnd vdd FILL
XFILL_26_DFFSR_115 gnd vdd FILL
XFILL_21_MUX2X1_2 gnd vdd FILL
XFILL_26_DFFSR_126 gnd vdd FILL
XFILL_26_DFFSR_137 gnd vdd FILL
XFILL_26_DFFSR_148 gnd vdd FILL
XFILL_26_DFFSR_159 gnd vdd FILL
XINVX1_102 INVX1_102/A gnd OAI22X1_7/A vdd INVX1
XINVX1_113 NOR2X1_13/Y gnd NOR2X1_24/B vdd INVX1
XFILL_5_NOR2X1_5 gnd vdd FILL
XINVX1_124 NOR2X1_24/Y gnd NOR2X1_35/B vdd INVX1
XINVX1_135 INVX1_135/A gnd NOR3X1_15/A vdd INVX1
XINVX1_146 INVX1_146/A gnd OAI21X1_4/A vdd INVX1
XINVX1_157 INVX1_157/A gnd INVX1_157/Y vdd INVX1
XFILL_15_MUX2X1_120 gnd vdd FILL
XINVX1_168 INVX1_168/A gnd INVX1_168/Y vdd INVX1
XINVX1_179 INVX1_179/A gnd INVX1_179/Y vdd INVX1
XFILL_29_DFFSR_50 gnd vdd FILL
XFILL_15_MUX2X1_131 gnd vdd FILL
XFILL_29_DFFSR_61 gnd vdd FILL
XFILL_17_INVX8_3 gnd vdd FILL
XFILL_15_MUX2X1_142 gnd vdd FILL
XFILL_29_DFFSR_72 gnd vdd FILL
XFILL_15_MUX2X1_153 gnd vdd FILL
XFILL_29_DFFSR_83 gnd vdd FILL
XFILL_22_NOR3X1_16 gnd vdd FILL
XFILL_15_MUX2X1_164 gnd vdd FILL
XFILL_22_NOR3X1_27 gnd vdd FILL
XFILL_29_DFFSR_94 gnd vdd FILL
XFILL_15_MUX2X1_175 gnd vdd FILL
XFILL_22_NOR3X1_38 gnd vdd FILL
XFILL_15_MUX2X1_186 gnd vdd FILL
XFILL_22_NOR3X1_49 gnd vdd FILL
XFILL_72_DFFSR_205 gnd vdd FILL
XFILL_72_DFFSR_216 gnd vdd FILL
XFILL_4_MUX2X1_3 gnd vdd FILL
XFILL_72_DFFSR_227 gnd vdd FILL
XFILL_49_1_0 gnd vdd FILL
XFILL_69_DFFSR_60 gnd vdd FILL
XFILL_72_DFFSR_238 gnd vdd FILL
XFILL_69_DFFSR_71 gnd vdd FILL
XFILL_69_DFFSR_82 gnd vdd FILL
XFILL_72_DFFSR_249 gnd vdd FILL
XFILL_21_DFFSR_5 gnd vdd FILL
XFILL_26_NOR3X1_15 gnd vdd FILL
XFILL_69_DFFSR_93 gnd vdd FILL
XFILL_26_NOR3X1_26 gnd vdd FILL
XFILL_26_NOR3X1_37 gnd vdd FILL
XFILL_26_NOR3X1_48 gnd vdd FILL
XFILL_76_DFFSR_204 gnd vdd FILL
XFILL_59_DFFSR_3 gnd vdd FILL
XFILL_76_DFFSR_215 gnd vdd FILL
XFILL_76_DFFSR_226 gnd vdd FILL
XFILL_76_DFFSR_237 gnd vdd FILL
XFILL_1_NOR3X1_9 gnd vdd FILL
XFILL_76_DFFSR_248 gnd vdd FILL
XFILL_11_DFFSR_170 gnd vdd FILL
XFILL_0_CLKBUF1_2 gnd vdd FILL
XFILL_76_DFFSR_259 gnd vdd FILL
XFILL_11_DFFSR_181 gnd vdd FILL
XFILL_34_4 gnd vdd FILL
XFILL_11_DFFSR_192 gnd vdd FILL
XFILL_38_DFFSR_70 gnd vdd FILL
XFILL_38_DFFSR_81 gnd vdd FILL
XFILL_38_DFFSR_92 gnd vdd FILL
XFILL_33_5_1 gnd vdd FILL
XFILL_27_3 gnd vdd FILL
XFILL_32_0_0 gnd vdd FILL
XFILL_4_CLKBUF1_1 gnd vdd FILL
XFILL_15_DFFSR_180 gnd vdd FILL
XFILL_15_DFFSR_191 gnd vdd FILL
XFILL_78_DFFSR_80 gnd vdd FILL
XFILL_78_DFFSR_91 gnd vdd FILL
XFILL_43_DFFSR_9 gnd vdd FILL
XFILL_5_MUX2X1_170 gnd vdd FILL
XFILL_5_MUX2X1_181 gnd vdd FILL
XFILL_5_MUX2X1_192 gnd vdd FILL
XFILL_19_DFFSR_190 gnd vdd FILL
XFILL_47_DFFSR_90 gnd vdd FILL
XFILL_61_DFFSR_270 gnd vdd FILL
XFILL_11_NAND2X1_14 gnd vdd FILL
XFILL_11_NAND2X1_25 gnd vdd FILL
XFILL_11_NAND2X1_36 gnd vdd FILL
XFILL_11_NAND2X1_47 gnd vdd FILL
XFILL_1_OAI21X1_6 gnd vdd FILL
XFILL_11_NAND2X1_58 gnd vdd FILL
XFILL_9_OAI22X1_19 gnd vdd FILL
XFILL_11_NAND2X1_69 gnd vdd FILL
XFILL_43_DFFSR_204 gnd vdd FILL
XFILL_43_DFFSR_215 gnd vdd FILL
XFILL_5_OAI21X1_5 gnd vdd FILL
XFILL_2_NOR2X1_30 gnd vdd FILL
XFILL_43_DFFSR_226 gnd vdd FILL
XFILL_2_NOR2X1_41 gnd vdd FILL
XFILL_2_NOR2X1_52 gnd vdd FILL
XFILL_43_DFFSR_237 gnd vdd FILL
XFILL_8_NAND3X1_40 gnd vdd FILL
XFILL_43_DFFSR_248 gnd vdd FILL
XFILL_2_NOR2X1_63 gnd vdd FILL
XFILL_8_NAND3X1_51 gnd vdd FILL
XFILL_8_NAND3X1_62 gnd vdd FILL
XFILL_2_NOR2X1_74 gnd vdd FILL
XFILL_24_5_1 gnd vdd FILL
XFILL_43_DFFSR_259 gnd vdd FILL
XFILL_8_NAND3X1_73 gnd vdd FILL
XFILL_2_NOR2X1_85 gnd vdd FILL
XFILL_70_DFFSR_104 gnd vdd FILL
XFILL_8_NAND3X1_84 gnd vdd FILL
XFILL_2_NOR2X1_96 gnd vdd FILL
XFILL_23_0_0 gnd vdd FILL
XFILL_8_NAND3X1_95 gnd vdd FILL
XFILL_47_DFFSR_203 gnd vdd FILL
XFILL_70_DFFSR_115 gnd vdd FILL
XFILL_5_BUFX4_8 gnd vdd FILL
XFILL_47_DFFSR_214 gnd vdd FILL
XFILL_9_OAI21X1_4 gnd vdd FILL
XFILL_70_DFFSR_126 gnd vdd FILL
XFILL_47_DFFSR_225 gnd vdd FILL
XFILL_70_DFFSR_137 gnd vdd FILL
XFILL_47_DFFSR_236 gnd vdd FILL
XFILL_6_NOR2X1_40 gnd vdd FILL
XFILL_10_OAI22X1_2 gnd vdd FILL
XFILL_70_DFFSR_148 gnd vdd FILL
XFILL_6_NOR2X1_51 gnd vdd FILL
XFILL_6_NOR2X1_62 gnd vdd FILL
XFILL_47_DFFSR_247 gnd vdd FILL
XFILL_70_DFFSR_159 gnd vdd FILL
XFILL_47_DFFSR_258 gnd vdd FILL
XFILL_6_NOR2X1_73 gnd vdd FILL
XFILL_47_DFFSR_269 gnd vdd FILL
XFILL_6_NOR2X1_84 gnd vdd FILL
XFILL_6_NOR2X1_95 gnd vdd FILL
XFILL_74_DFFSR_103 gnd vdd FILL
XFILL_74_DFFSR_114 gnd vdd FILL
XFILL_74_DFFSR_125 gnd vdd FILL
XFILL_74_DFFSR_136 gnd vdd FILL
XFILL_15_AOI21X1_14 gnd vdd FILL
XFILL_14_OAI22X1_1 gnd vdd FILL
XFILL_74_DFFSR_147 gnd vdd FILL
XFILL_74_DFFSR_158 gnd vdd FILL
XFILL_15_AOI21X1_25 gnd vdd FILL
XFILL_74_DFFSR_169 gnd vdd FILL
XFILL_1_NAND2X1_20 gnd vdd FILL
XFILL_15_AOI21X1_36 gnd vdd FILL
XFILL_1_NAND2X1_31 gnd vdd FILL
XFILL_15_AOI21X1_47 gnd vdd FILL
XFILL_78_DFFSR_102 gnd vdd FILL
XFILL_1_NAND2X1_42 gnd vdd FILL
XFILL_15_AOI21X1_58 gnd vdd FILL
XFILL_15_AOI21X1_69 gnd vdd FILL
XFILL_1_NAND2X1_53 gnd vdd FILL
XFILL_78_DFFSR_113 gnd vdd FILL
XFILL_78_DFFSR_124 gnd vdd FILL
XFILL_12_BUFX4_16 gnd vdd FILL
XFILL_1_NAND2X1_64 gnd vdd FILL
XFILL_12_BUFX4_27 gnd vdd FILL
XFILL_1_NAND2X1_75 gnd vdd FILL
XFILL_78_DFFSR_135 gnd vdd FILL
XFILL_1_NAND2X1_86 gnd vdd FILL
XFILL_78_DFFSR_146 gnd vdd FILL
XFILL_12_BUFX4_38 gnd vdd FILL
XFILL_78_DFFSR_157 gnd vdd FILL
XFILL_12_BUFX4_49 gnd vdd FILL
XFILL_78_DFFSR_168 gnd vdd FILL
XFILL_78_DFFSR_179 gnd vdd FILL
XFILL_1_BUFX2_4 gnd vdd FILL
XFILL_7_6_1 gnd vdd FILL
XFILL_6_1_0 gnd vdd FILL
XFILL_6_NAND3X1_110 gnd vdd FILL
XFILL_6_NAND3X1_121 gnd vdd FILL
XFILL_6_NAND3X1_132 gnd vdd FILL
XFILL_2_NAND2X1_7 gnd vdd FILL
XFILL_60_DFFSR_3 gnd vdd FILL
XFILL_27_CLKBUF1_30 gnd vdd FILL
XFILL_27_CLKBUF1_41 gnd vdd FILL
XFILL_6_INVX1_17 gnd vdd FILL
XFILL_6_NAND2X1_6 gnd vdd FILL
XFILL_6_INVX1_28 gnd vdd FILL
XFILL_10_DFFSR_204 gnd vdd FILL
XFILL_10_DFFSR_215 gnd vdd FILL
XFILL_15_5_1 gnd vdd FILL
XFILL_6_INVX1_39 gnd vdd FILL
XFILL_18_MUX2X1_108 gnd vdd FILL
XFILL_18_MUX2X1_119 gnd vdd FILL
XFILL_5_AOI21X1_20 gnd vdd FILL
XFILL_2_MUX2X1_70 gnd vdd FILL
XFILL_5_AOI21X1_31 gnd vdd FILL
XFILL_10_DFFSR_226 gnd vdd FILL
XFILL_10_DFFSR_237 gnd vdd FILL
XFILL_14_0_0 gnd vdd FILL
XFILL_2_MUX2X1_81 gnd vdd FILL
XFILL_5_AOI21X1_42 gnd vdd FILL
XFILL_10_DFFSR_248 gnd vdd FILL
XFILL_2_MUX2X1_92 gnd vdd FILL
XFILL_15_OAI22X1_11 gnd vdd FILL
XFILL_5_AOI21X1_53 gnd vdd FILL
XFILL_10_DFFSR_259 gnd vdd FILL
XFILL_5_AOI21X1_64 gnd vdd FILL
XFILL_5_AOI21X1_75 gnd vdd FILL
XFILL_15_OAI22X1_22 gnd vdd FILL
XFILL_63_DFFSR_190 gnd vdd FILL
XFILL_15_OAI22X1_33 gnd vdd FILL
XFILL_15_OAI22X1_44 gnd vdd FILL
XFILL_14_DFFSR_203 gnd vdd FILL
XFILL_11_NAND3X1_3 gnd vdd FILL
XFILL_14_DFFSR_214 gnd vdd FILL
XFILL_14_DFFSR_225 gnd vdd FILL
XFILL_6_MUX2X1_80 gnd vdd FILL
XFILL_14_DFFSR_236 gnd vdd FILL
XFILL_8_NOR2X1_130 gnd vdd FILL
XFILL_8_NOR2X1_141 gnd vdd FILL
XFILL_14_DFFSR_247 gnd vdd FILL
XFILL_6_MUX2X1_91 gnd vdd FILL
XDFFSR_108 INVX1_189/A DFFSR_78/CLK DFFSR_78/R vdd DFFSR_108/D gnd vdd DFFSR
XFILL_25_DFFSR_6 gnd vdd FILL
XFILL_14_DFFSR_258 gnd vdd FILL
XFILL_8_NOR2X1_152 gnd vdd FILL
XFILL_14_DFFSR_269 gnd vdd FILL
XDFFSR_119 INVX1_181/A DFFSR_52/CLK DFFSR_56/R vdd DFFSR_119/D gnd vdd DFFSR
XFILL_4_BUFX4_15 gnd vdd FILL
XFILL_8_NOR2X1_163 gnd vdd FILL
XFILL_8_NOR2X1_174 gnd vdd FILL
XFILL_4_BUFX4_26 gnd vdd FILL
XFILL_82_DFFSR_7 gnd vdd FILL
XFILL_41_DFFSR_103 gnd vdd FILL
XFILL_4_BUFX4_37 gnd vdd FILL
XFILL_18_DFFSR_202 gnd vdd FILL
XFILL_4_BUFX4_48 gnd vdd FILL
XFILL_15_NAND3X1_2 gnd vdd FILL
XFILL_8_NOR2X1_185 gnd vdd FILL
XFILL_18_DFFSR_213 gnd vdd FILL
XFILL_41_DFFSR_114 gnd vdd FILL
XFILL_8_NOR2X1_196 gnd vdd FILL
XFILL_4_BUFX4_59 gnd vdd FILL
XFILL_18_DFFSR_224 gnd vdd FILL
XFILL_1_INVX2_4 gnd vdd FILL
XFILL_41_DFFSR_125 gnd vdd FILL
XFILL_41_DFFSR_136 gnd vdd FILL
XFILL_18_DFFSR_235 gnd vdd FILL
XFILL_41_DFFSR_147 gnd vdd FILL
XFILL_41_DFFSR_158 gnd vdd FILL
XFILL_18_DFFSR_246 gnd vdd FILL
XFILL_18_DFFSR_257 gnd vdd FILL
XFILL_18_DFFSR_268 gnd vdd FILL
XFILL_41_DFFSR_169 gnd vdd FILL
XFILL_45_DFFSR_102 gnd vdd FILL
XFILL_45_DFFSR_113 gnd vdd FILL
XFILL_45_DFFSR_124 gnd vdd FILL
XFILL_45_DFFSR_135 gnd vdd FILL
XFILL_45_DFFSR_146 gnd vdd FILL
XFILL_45_DFFSR_157 gnd vdd FILL
XFILL_45_DFFSR_168 gnd vdd FILL
XFILL_45_DFFSR_179 gnd vdd FILL
XFILL_8_MUX2X1_103 gnd vdd FILL
XFILL_49_DFFSR_101 gnd vdd FILL
XFILL_8_MUX2X1_114 gnd vdd FILL
XFILL_49_DFFSR_112 gnd vdd FILL
XFILL_8_MUX2X1_125 gnd vdd FILL
XFILL_49_DFFSR_123 gnd vdd FILL
XFILL_8_MUX2X1_136 gnd vdd FILL
XFILL_49_DFFSR_134 gnd vdd FILL
XFILL_49_DFFSR_145 gnd vdd FILL
XFILL_11_AND2X2_3 gnd vdd FILL
XFILL_8_MUX2X1_147 gnd vdd FILL
XFILL_49_DFFSR_156 gnd vdd FILL
XFILL_8_MUX2X1_158 gnd vdd FILL
XFILL_11_AOI22X1_8 gnd vdd FILL
XNOR3X1_19 INVX1_39/Y NOR3X1_29/B NOR3X1_6/C gnd NOR3X1_20/A vdd NOR3X1
XFILL_49_DFFSR_167 gnd vdd FILL
XFILL_8_MUX2X1_169 gnd vdd FILL
XFILL_49_DFFSR_178 gnd vdd FILL
XFILL_65_4_1 gnd vdd FILL
XFILL_5_OAI22X1_50 gnd vdd FILL
XFILL_49_DFFSR_189 gnd vdd FILL
XFILL_9_OAI21X1_30 gnd vdd FILL
XFILL_9_OAI21X1_41 gnd vdd FILL
XFILL_15_AOI22X1_7 gnd vdd FILL
XFILL_32_1 gnd vdd FILL
XFILL_19_AOI22X1_6 gnd vdd FILL
XFILL_30_DFFSR_190 gnd vdd FILL
XFILL_39_DFFSR_15 gnd vdd FILL
XFILL_39_DFFSR_26 gnd vdd FILL
XFILL_39_DFFSR_37 gnd vdd FILL
XFILL_39_DFFSR_48 gnd vdd FILL
XFILL_39_DFFSR_59 gnd vdd FILL
XFILL_79_DFFSR_14 gnd vdd FILL
XFILL_79_DFFSR_25 gnd vdd FILL
XFILL_79_DFFSR_36 gnd vdd FILL
XFILL_79_DFFSR_47 gnd vdd FILL
XFILL_79_DFFSR_58 gnd vdd FILL
XFILL_79_DFFSR_69 gnd vdd FILL
XFILL_2_INVX1_10 gnd vdd FILL
XFILL_2_INVX1_21 gnd vdd FILL
XFILL_12_DFFSR_102 gnd vdd FILL
XFILL_2_INVX1_32 gnd vdd FILL
XFILL_2_INVX1_43 gnd vdd FILL
XFILL_12_DFFSR_113 gnd vdd FILL
XFILL_3_AND2X2_2 gnd vdd FILL
XFILL_9_BUFX4_9 gnd vdd FILL
XFILL_2_INVX1_54 gnd vdd FILL
XFILL_12_DFFSR_124 gnd vdd FILL
XFILL_2_INVX1_65 gnd vdd FILL
XFILL_12_DFFSR_135 gnd vdd FILL
XFILL_2_INVX1_76 gnd vdd FILL
XFILL_12_DFFSR_146 gnd vdd FILL
XFILL_48_DFFSR_13 gnd vdd FILL
XFILL_12_DFFSR_157 gnd vdd FILL
XFILL_48_DFFSR_24 gnd vdd FILL
XFILL_2_INVX1_87 gnd vdd FILL
XFILL_48_DFFSR_35 gnd vdd FILL
XFILL_2_INVX1_98 gnd vdd FILL
XFILL_48_DFFSR_46 gnd vdd FILL
XFILL_12_DFFSR_168 gnd vdd FILL
XFILL_12_DFFSR_179 gnd vdd FILL
XFILL_16_DFFSR_101 gnd vdd FILL
XFILL_48_DFFSR_57 gnd vdd FILL
XFILL_48_DFFSR_68 gnd vdd FILL
XFILL_16_DFFSR_112 gnd vdd FILL
XFILL_48_DFFSR_79 gnd vdd FILL
XFILL_0_NAND3X1_17 gnd vdd FILL
XFILL_16_DFFSR_123 gnd vdd FILL
XFILL_16_DFFSR_134 gnd vdd FILL
XFILL_56_4_1 gnd vdd FILL
XFILL_0_NAND3X1_28 gnd vdd FILL
XFILL_16_DFFSR_145 gnd vdd FILL
XFILL_0_NAND3X1_39 gnd vdd FILL
XFILL_16_DFFSR_156 gnd vdd FILL
XFILL_16_DFFSR_167 gnd vdd FILL
XFILL_0_BUFX4_30 gnd vdd FILL
XFILL_4_NAND2X1_19 gnd vdd FILL
XFILL_16_DFFSR_178 gnd vdd FILL
XFILL_0_BUFX4_41 gnd vdd FILL
XFILL_17_DFFSR_12 gnd vdd FILL
XFILL_0_BUFX4_52 gnd vdd FILL
XFILL_16_DFFSR_189 gnd vdd FILL
XFILL_0_BUFX4_63 gnd vdd FILL
XFILL_17_DFFSR_23 gnd vdd FILL
XFILL_17_DFFSR_34 gnd vdd FILL
XFILL_0_BUFX4_74 gnd vdd FILL
XFILL_17_DFFSR_45 gnd vdd FILL
XFILL_17_DFFSR_56 gnd vdd FILL
XFILL_0_BUFX4_85 gnd vdd FILL
XFILL_0_BUFX4_96 gnd vdd FILL
XFILL_17_DFFSR_67 gnd vdd FILL
XFILL_1_BUFX4_105 gnd vdd FILL
XFILL_17_DFFSR_78 gnd vdd FILL
XFILL_17_DFFSR_89 gnd vdd FILL
XFILL_14_MUX2X1_150 gnd vdd FILL
XFILL_14_MUX2X1_161 gnd vdd FILL
XFILL_9_CLKBUF1_9 gnd vdd FILL
XFILL_12_NOR3X1_13 gnd vdd FILL
XFILL_57_DFFSR_11 gnd vdd FILL
XFILL_12_NOR3X1_24 gnd vdd FILL
XFILL_14_MUX2X1_172 gnd vdd FILL
XFILL_5_BUFX2_5 gnd vdd FILL
XFILL_12_NOR3X1_35 gnd vdd FILL
XFILL_57_DFFSR_22 gnd vdd FILL
XFILL_57_DFFSR_33 gnd vdd FILL
XFILL_14_MUX2X1_183 gnd vdd FILL
XFILL_62_DFFSR_202 gnd vdd FILL
XFILL_28_NOR3X1_8 gnd vdd FILL
XFILL_12_NOR3X1_46 gnd vdd FILL
XFILL_14_MUX2X1_194 gnd vdd FILL
XFILL_57_DFFSR_44 gnd vdd FILL
XFILL_57_DFFSR_55 gnd vdd FILL
XFILL_62_DFFSR_213 gnd vdd FILL
XFILL_57_DFFSR_66 gnd vdd FILL
XFILL_62_DFFSR_224 gnd vdd FILL
XFILL_62_DFFSR_235 gnd vdd FILL
XFILL_5_BUFX4_104 gnd vdd FILL
XFILL_57_DFFSR_77 gnd vdd FILL
XFILL_57_DFFSR_88 gnd vdd FILL
XFILL_62_DFFSR_246 gnd vdd FILL
XFILL_57_DFFSR_99 gnd vdd FILL
XFILL_16_NOR3X1_12 gnd vdd FILL
XFILL_62_DFFSR_257 gnd vdd FILL
XFILL_62_DFFSR_268 gnd vdd FILL
XFILL_16_NOR3X1_23 gnd vdd FILL
XFILL_16_NOR3X1_34 gnd vdd FILL
XFILL_16_NOR3X1_45 gnd vdd FILL
XFILL_66_DFFSR_201 gnd vdd FILL
XFILL_64_DFFSR_4 gnd vdd FILL
XFILL_2_NOR2X1_9 gnd vdd FILL
XFILL_66_DFFSR_212 gnd vdd FILL
XFILL_26_DFFSR_10 gnd vdd FILL
XFILL_26_DFFSR_21 gnd vdd FILL
XFILL_66_DFFSR_223 gnd vdd FILL
XFILL_66_DFFSR_234 gnd vdd FILL
XFILL_9_BUFX4_103 gnd vdd FILL
XFILL_26_DFFSR_32 gnd vdd FILL
XFILL_26_DFFSR_43 gnd vdd FILL
XFILL_3_OR2X2_1 gnd vdd FILL
XFILL_66_DFFSR_245 gnd vdd FILL
XFILL_66_DFFSR_256 gnd vdd FILL
XFILL_26_DFFSR_54 gnd vdd FILL
XFILL_66_DFFSR_267 gnd vdd FILL
XFILL_26_DFFSR_65 gnd vdd FILL
XFILL_26_DFFSR_76 gnd vdd FILL
XFILL_21_CLKBUF1_8 gnd vdd FILL
XFILL_26_DFFSR_87 gnd vdd FILL
XFILL_26_DFFSR_98 gnd vdd FILL
XFILL_8_AOI21X1_19 gnd vdd FILL
XFILL_66_DFFSR_20 gnd vdd FILL
XFILL_66_DFFSR_31 gnd vdd FILL
XFILL_66_DFFSR_42 gnd vdd FILL
XFILL_1_MUX2X1_7 gnd vdd FILL
XFILL_66_DFFSR_53 gnd vdd FILL
XFILL_66_DFFSR_64 gnd vdd FILL
XFILL_25_CLKBUF1_7 gnd vdd FILL
XFILL_66_DFFSR_75 gnd vdd FILL
XFILL_66_DFFSR_86 gnd vdd FILL
XFILL_3_NOR2X1_17 gnd vdd FILL
XNAND3X1_30 OAI21X1_41/A AND2X2_7/Y NAND3X1_30/C gnd AOI22X1_2/C vdd NAND3X1
XFILL_66_DFFSR_97 gnd vdd FILL
XFILL_3_NOR2X1_28 gnd vdd FILL
XNAND3X1_41 DFFSR_19/Q BUFX4_8/Y NOR2X1_34/Y gnd NAND3X1_46/B vdd NAND3X1
XFILL_9_DFFSR_11 gnd vdd FILL
XFILL_3_NOR2X1_39 gnd vdd FILL
XNAND3X1_52 AND2X2_6/B AND2X2_6/A BUFX4_6/Y gnd INVX1_121/A vdd NAND3X1
XFILL_9_DFFSR_22 gnd vdd FILL
XFILL_7_NAND3X1_100 gnd vdd FILL
XFILL_29_DFFSR_7 gnd vdd FILL
XNAND3X1_63 BUFX4_58/Y AND2X2_3/B NAND3X1_2/C gnd OAI22X1_3/D vdd NAND3X1
XNAND3X1_74 DFFSR_81/Q BUFX4_1/Y NOR2X1_44/Y gnd OAI21X1_5/C vdd NAND3X1
XFILL_9_DFFSR_33 gnd vdd FILL
XFILL_7_NAND3X1_111 gnd vdd FILL
XFILL_47_4_1 gnd vdd FILL
XFILL_86_DFFSR_8 gnd vdd FILL
XNAND3X1_85 AOI22X1_7/Y NAND3X1_85/B NOR3X1_17/Y gnd NOR3X1_18/A vdd NAND3X1
XFILL_7_NAND3X1_122 gnd vdd FILL
XFILL_9_DFFSR_44 gnd vdd FILL
XFILL_9_DFFSR_55 gnd vdd FILL
XNAND3X1_96 DFFSR_104/Q BUFX4_2/Y NOR2X1_29/Y gnd OAI21X1_17/C vdd NAND3X1
XFILL_35_DFFSR_30 gnd vdd FILL
XFILL_29_CLKBUF1_6 gnd vdd FILL
XFILL_9_DFFSR_66 gnd vdd FILL
XFILL_35_DFFSR_41 gnd vdd FILL
XFILL_9_DFFSR_77 gnd vdd FILL
XNOR2X1_30 NOR3X1_2/C NOR2X1_37/B gnd NOR2X1_30/Y vdd NOR2X1
XFILL_7_NOR2X1_16 gnd vdd FILL
XNOR2X1_41 NOR3X1_49/B NOR2X1_41/B gnd NOR2X1_41/Y vdd NOR2X1
XFILL_7_NOR2X1_27 gnd vdd FILL
XFILL_35_DFFSR_52 gnd vdd FILL
XFILL_5_INVX2_5 gnd vdd FILL
XFILL_35_DFFSR_63 gnd vdd FILL
XFILL_9_DFFSR_88 gnd vdd FILL
XNOR2X1_52 NOR3X1_6/C NOR2X1_52/B gnd NOR2X1_52/Y vdd NOR2X1
XFILL_9_DFFSR_99 gnd vdd FILL
XFILL_35_DFFSR_74 gnd vdd FILL
XFILL_7_NOR2X1_38 gnd vdd FILL
XFILL_35_DFFSR_85 gnd vdd FILL
XNOR2X1_63 NOR2X1_63/A OAI22X1_9/Y gnd NOR2X1_63/Y vdd NOR2X1
XFILL_7_NOR2X1_49 gnd vdd FILL
XNOR2X1_74 NOR2X1_74/A NOR2X1_74/B gnd NOR2X1_74/Y vdd NOR2X1
XFILL_35_DFFSR_96 gnd vdd FILL
XNOR2X1_85 NOR2X1_85/A NOR2X1_85/B gnd NOR2X1_85/Y vdd NOR2X1
XNOR2X1_96 NOR2X1_96/A NOR2X1_96/B gnd NOR2X1_96/Y vdd NOR2X1
XFILL_75_DFFSR_40 gnd vdd FILL
XFILL_75_DFFSR_51 gnd vdd FILL
XFILL_0_NOR2X1_107 gnd vdd FILL
XFILL_0_NOR2X1_118 gnd vdd FILL
XFILL_75_DFFSR_62 gnd vdd FILL
XFILL_0_NOR2X1_129 gnd vdd FILL
XFILL_75_DFFSR_73 gnd vdd FILL
XFILL_75_DFFSR_84 gnd vdd FILL
XFILL_75_DFFSR_95 gnd vdd FILL
XFILL_3_INVX1_3 gnd vdd FILL
XFILL_10_NAND2X1_11 gnd vdd FILL
XFILL_30_3_1 gnd vdd FILL
XFILL_10_NAND2X1_22 gnd vdd FILL
XFILL_10_NAND2X1_33 gnd vdd FILL
XFILL_10_NAND2X1_44 gnd vdd FILL
XFILL_10_NAND2X1_55 gnd vdd FILL
XFILL_10_NAND2X1_66 gnd vdd FILL
XFILL_15_NOR3X1_3 gnd vdd FILL
XFILL_19_OAI22X1_9 gnd vdd FILL
XFILL_8_OAI22X1_16 gnd vdd FILL
XFILL_44_DFFSR_50 gnd vdd FILL
XFILL_10_NAND2X1_77 gnd vdd FILL
XFILL_8_OAI22X1_27 gnd vdd FILL
XFILL_44_DFFSR_61 gnd vdd FILL
XFILL_10_NAND2X1_88 gnd vdd FILL
XFILL_8_OAI22X1_38 gnd vdd FILL
XFILL_44_DFFSR_72 gnd vdd FILL
XFILL_44_DFFSR_83 gnd vdd FILL
XFILL_8_OAI22X1_49 gnd vdd FILL
XFILL_44_DFFSR_94 gnd vdd FILL
XFILL_33_DFFSR_201 gnd vdd FILL
XFILL_33_DFFSR_212 gnd vdd FILL
XFILL_33_DFFSR_223 gnd vdd FILL
XFILL_33_DFFSR_234 gnd vdd FILL
XFILL_33_DFFSR_245 gnd vdd FILL
XFILL_84_DFFSR_60 gnd vdd FILL
XFILL_33_DFFSR_256 gnd vdd FILL
XFILL_84_DFFSR_71 gnd vdd FILL
XFILL_33_DFFSR_267 gnd vdd FILL
XFILL_7_NAND3X1_70 gnd vdd FILL
XFILL_84_DFFSR_82 gnd vdd FILL
XFILL_60_DFFSR_101 gnd vdd FILL
XFILL_84_DFFSR_93 gnd vdd FILL
XFILL_7_NAND3X1_81 gnd vdd FILL
XFILL_7_NAND3X1_92 gnd vdd FILL
XFILL_37_DFFSR_200 gnd vdd FILL
XFILL_13_DFFSR_60 gnd vdd FILL
XFILL_60_DFFSR_112 gnd vdd FILL
XFILL_37_DFFSR_211 gnd vdd FILL
XFILL_13_DFFSR_71 gnd vdd FILL
XFILL_37_DFFSR_222 gnd vdd FILL
XFILL_60_DFFSR_123 gnd vdd FILL
XFILL_13_DFFSR_82 gnd vdd FILL
XFILL_60_DFFSR_134 gnd vdd FILL
XFILL_37_DFFSR_233 gnd vdd FILL
XFILL_13_DFFSR_93 gnd vdd FILL
XFILL_60_DFFSR_145 gnd vdd FILL
XFILL_37_DFFSR_244 gnd vdd FILL
XFILL_60_DFFSR_156 gnd vdd FILL
XFILL_37_DFFSR_255 gnd vdd FILL
XFILL_60_DFFSR_167 gnd vdd FILL
XFILL_3_MUX2X1_13 gnd vdd FILL
XFILL_24_NOR3X1_1 gnd vdd FILL
XFILL_37_DFFSR_266 gnd vdd FILL
XNAND2X1_7 INVX2_1/A INVX1_2/A gnd NAND2X1_7/Y vdd NAND2X1
XFILL_60_DFFSR_178 gnd vdd FILL
XFILL_3_MUX2X1_24 gnd vdd FILL
XFILL_1_OAI21X1_18 gnd vdd FILL
XFILL_64_DFFSR_100 gnd vdd FILL
XFILL_60_DFFSR_189 gnd vdd FILL
XFILL_1_OAI21X1_29 gnd vdd FILL
XFILL_3_MUX2X1_35 gnd vdd FILL
XFILL_64_DFFSR_111 gnd vdd FILL
XFILL_19_CLKBUF1_14 gnd vdd FILL
XFILL_19_CLKBUF1_25 gnd vdd FILL
XFILL_53_DFFSR_70 gnd vdd FILL
XFILL_64_DFFSR_122 gnd vdd FILL
XFILL_3_MUX2X1_46 gnd vdd FILL
XFILL_38_4_1 gnd vdd FILL
XFILL_53_DFFSR_81 gnd vdd FILL
XFILL_3_MUX2X1_57 gnd vdd FILL
XFILL_19_CLKBUF1_36 gnd vdd FILL
XFILL_64_DFFSR_133 gnd vdd FILL
XFILL_3_MUX2X1_68 gnd vdd FILL
XFILL_14_AOI21X1_11 gnd vdd FILL
XFILL_53_DFFSR_92 gnd vdd FILL
XFILL_64_DFFSR_144 gnd vdd FILL
XFILL_3_MUX2X1_79 gnd vdd FILL
XFILL_64_DFFSR_155 gnd vdd FILL
XFILL_14_AOI21X1_22 gnd vdd FILL
XFILL_64_DFFSR_166 gnd vdd FILL
XFILL_14_AOI21X1_33 gnd vdd FILL
XFILL_7_MUX2X1_12 gnd vdd FILL
XFILL_14_AOI21X1_44 gnd vdd FILL
XFILL_7_MUX2X1_23 gnd vdd FILL
XFILL_64_DFFSR_177 gnd vdd FILL
XFILL_64_DFFSR_188 gnd vdd FILL
XFILL_14_AOI21X1_55 gnd vdd FILL
XFILL_14_AOI21X1_66 gnd vdd FILL
XFILL_0_NAND2X1_50 gnd vdd FILL
XFILL_7_MUX2X1_34 gnd vdd FILL
XNOR2X1_120 INVX1_139/A NOR2X1_21/A gnd INVX4_1/A vdd NOR2X1
XFILL_68_DFFSR_110 gnd vdd FILL
XFILL_64_DFFSR_199 gnd vdd FILL
XFILL_7_MUX2X1_45 gnd vdd FILL
XFILL_68_DFFSR_121 gnd vdd FILL
XFILL_0_NAND2X1_61 gnd vdd FILL
XFILL_68_DFFSR_132 gnd vdd FILL
XMUX2X1_70 INVX1_83/Y BUFX4_75/Y MUX2X1_71/S gnd MUX2X1_70/Y vdd MUX2X1
XFILL_0_NAND2X1_72 gnd vdd FILL
XFILL_14_AOI21X1_77 gnd vdd FILL
XFILL_7_MUX2X1_56 gnd vdd FILL
XNOR2X1_131 DFFSR_139/Q AOI21X1_7/B gnd AOI21X1_4/C vdd NOR2X1
XMUX2X1_81 BUFX4_64/Y INVX1_94/Y NOR2X1_28/B gnd MUX2X1_81/Y vdd MUX2X1
XFILL_0_NAND2X1_83 gnd vdd FILL
XFILL_7_MUX2X1_67 gnd vdd FILL
XNOR2X1_142 NAND2X1_3/Y INVX1_174/Y gnd NOR2X1_142/Y vdd NOR2X1
XFILL_68_DFFSR_143 gnd vdd FILL
XMUX2X1_92 MUX2X1_92/A BUFX4_86/Y MUX2X1_95/S gnd MUX2X1_92/Y vdd MUX2X1
XFILL_7_MUX2X1_78 gnd vdd FILL
XNOR2X1_153 DFFSR_102/Q NOR2X1_153/B gnd NOR2X1_153/Y vdd NOR2X1
XFILL_0_NAND2X1_94 gnd vdd FILL
XFILL_68_DFFSR_154 gnd vdd FILL
XNOR2X1_164 NOR2X1_25/A NAND2X1_3/Y gnd NOR2X1_164/Y vdd NOR2X1
XFILL_68_DFFSR_165 gnd vdd FILL
XFILL_7_MUX2X1_89 gnd vdd FILL
XFILL_22_DFFSR_80 gnd vdd FILL
XNOR2X1_175 NOR2X1_7/B INVX1_2/Y gnd MUX2X1_14/S vdd NOR2X1
XFILL_68_DFFSR_176 gnd vdd FILL
XFILL_22_DFFSR_91 gnd vdd FILL
XNOR2X1_186 NOR2X1_57/A NOR2X1_7/B gnd NOR2X1_190/B vdd NOR2X1
XNOR2X1_197 NOR2X1_7/B INVX1_205/Y gnd MUX2X1_20/S vdd NOR2X1
XFILL_7_NOR3X1_2 gnd vdd FILL
XFILL_68_DFFSR_187 gnd vdd FILL
XFILL_68_DFFSR_198 gnd vdd FILL
XFILL_21_3_1 gnd vdd FILL
XFILL_62_DFFSR_90 gnd vdd FILL
XFILL_46_DFFSR_1 gnd vdd FILL
XMUX2X1_104 NOR3X1_46/A BUFX4_98/Y NAND2X1_16/Y gnd DFFSR_46/D vdd MUX2X1
XMUX2X1_115 BUFX4_76/Y INVX1_157/Y NOR2X1_128/Y gnd DFFSR_145/D vdd MUX2X1
XFILL_5_DFFSR_70 gnd vdd FILL
XFILL_9_CLKBUF1_20 gnd vdd FILL
XFILL_23_MUX2X1_10 gnd vdd FILL
XMUX2X1_126 INVX1_170/Y MUX2X1_4/B NAND2X1_89/Y gnd DFFSR_126/D vdd MUX2X1
XFILL_5_DFFSR_81 gnd vdd FILL
XFILL_23_MUX2X1_21 gnd vdd FILL
XFILL_5_DFFSR_92 gnd vdd FILL
XFILL_9_CLKBUF1_31 gnd vdd FILL
XFILL_9_CLKBUF1_42 gnd vdd FILL
XMUX2X1_137 BUFX4_72/Y INVX1_181/Y NOR2X1_139/Y gnd DFFSR_119/D vdd MUX2X1
XMUX2X1_148 BUFX4_81/Y OAI21X1_6/A NOR2X1_154/Y gnd DFFSR_94/D vdd MUX2X1
XFILL_23_MUX2X1_32 gnd vdd FILL
XFILL_17_MUX2X1_105 gnd vdd FILL
XFILL_17_MUX2X1_116 gnd vdd FILL
XMUX2X1_159 BUFX4_78/Y INVX1_203/Y NOR2X1_156/Y gnd DFFSR_87/D vdd MUX2X1
XFILL_23_MUX2X1_43 gnd vdd FILL
XFILL_23_MUX2X1_54 gnd vdd FILL
XFILL_17_MUX2X1_127 gnd vdd FILL
XFILL_23_MUX2X1_65 gnd vdd FILL
XFILL_23_MUX2X1_76 gnd vdd FILL
XFILL_17_MUX2X1_138 gnd vdd FILL
XFILL_17_MUX2X1_149 gnd vdd FILL
XFILL_4_AOI21X1_50 gnd vdd FILL
XFILL_23_MUX2X1_87 gnd vdd FILL
XFILL_4_AOI21X1_61 gnd vdd FILL
XFILL_9_BUFX2_6 gnd vdd FILL
XFILL_4_AOI21X1_72 gnd vdd FILL
XFILL_23_MUX2X1_98 gnd vdd FILL
XFILL_14_OAI22X1_30 gnd vdd FILL
XFILL_14_OAI22X1_41 gnd vdd FILL
XINVX1_11 INVX1_11/A gnd INVX1_11/Y vdd INVX1
XINVX1_22 INVX1_22/A gnd MUX2X1_9/B vdd INVX1
XINVX1_33 INVX1_33/A gnd INVX1_33/Y vdd INVX1
XINVX1_44 INVX1_44/A gnd INVX1_44/Y vdd INVX1
XINVX1_55 INVX1_55/A gnd INVX1_55/Y vdd INVX1
XFILL_30_DFFSR_7 gnd vdd FILL
XINVX1_66 INVX1_66/A gnd INVX1_66/Y vdd INVX1
XFILL_7_NOR2X1_160 gnd vdd FILL
XINVX1_77 INVX1_77/A gnd INVX1_77/Y vdd INVX1
XINVX1_88 INVX1_88/A gnd INVX1_88/Y vdd INVX1
XFILL_7_NOR2X1_171 gnd vdd FILL
XFILL_29_4_1 gnd vdd FILL
XINVX1_99 INVX1_99/A gnd INVX1_99/Y vdd INVX1
XFILL_31_DFFSR_100 gnd vdd FILL
XFILL_4_4_1 gnd vdd FILL
XFILL_7_NOR2X1_182 gnd vdd FILL
XFILL_31_DFFSR_111 gnd vdd FILL
XFILL_68_DFFSR_5 gnd vdd FILL
XFILL_7_NOR2X1_193 gnd vdd FILL
XFILL_31_DFFSR_122 gnd vdd FILL
XFILL_31_DFFSR_133 gnd vdd FILL
XFILL_31_DFFSR_144 gnd vdd FILL
XFILL_31_DFFSR_155 gnd vdd FILL
XFILL_31_DFFSR_166 gnd vdd FILL
XFILL_31_DFFSR_177 gnd vdd FILL
XFILL_0_DFFSR_190 gnd vdd FILL
XFILL_31_DFFSR_188 gnd vdd FILL
XFILL_35_DFFSR_110 gnd vdd FILL
XFILL_31_DFFSR_199 gnd vdd FILL
XFILL_35_DFFSR_121 gnd vdd FILL
XFILL_35_DFFSR_132 gnd vdd FILL
XFILL_35_DFFSR_143 gnd vdd FILL
XFILL_35_DFFSR_154 gnd vdd FILL
XFILL_35_DFFSR_165 gnd vdd FILL
XFILL_35_DFFSR_176 gnd vdd FILL
XFILL_12_3_1 gnd vdd FILL
XFILL_7_MUX2X1_100 gnd vdd FILL
XFILL_35_DFFSR_187 gnd vdd FILL
XFILL_7_MUX2X1_111 gnd vdd FILL
XFILL_35_DFFSR_198 gnd vdd FILL
XFILL_7_MUX2X1_122 gnd vdd FILL
XFILL_39_DFFSR_120 gnd vdd FILL
XFILL_1_BUFX4_19 gnd vdd FILL
XFILL_39_DFFSR_131 gnd vdd FILL
XFILL_7_MUX2X1_133 gnd vdd FILL
XFILL_7_MUX2X1_144 gnd vdd FILL
XFILL_39_DFFSR_142 gnd vdd FILL
XFILL_7_MUX2X1_155 gnd vdd FILL
XFILL_39_DFFSR_153 gnd vdd FILL
XFILL_7_MUX2X1_166 gnd vdd FILL
XFILL_39_DFFSR_164 gnd vdd FILL
XFILL_39_DFFSR_175 gnd vdd FILL
XFILL_7_MUX2X1_177 gnd vdd FILL
XFILL_31_NOR3X1_11 gnd vdd FILL
XFILL_39_DFFSR_186 gnd vdd FILL
XFILL_7_MUX2X1_188 gnd vdd FILL
XFILL_31_NOR3X1_22 gnd vdd FILL
XFILL_39_DFFSR_197 gnd vdd FILL
XFILL_31_NOR3X1_33 gnd vdd FILL
XFILL_31_NOR3X1_44 gnd vdd FILL
XFILL_81_DFFSR_200 gnd vdd FILL
XFILL_81_DFFSR_211 gnd vdd FILL
XFILL_81_DFFSR_222 gnd vdd FILL
XFILL_81_DFFSR_233 gnd vdd FILL
XFILL_81_DFFSR_244 gnd vdd FILL
XFILL_81_DFFSR_255 gnd vdd FILL
XFILL_81_DFFSR_266 gnd vdd FILL
XFILL_85_DFFSR_210 gnd vdd FILL
XFILL_85_DFFSR_221 gnd vdd FILL
XFILL_12_AOI21X1_6 gnd vdd FILL
XFILL_85_DFFSR_232 gnd vdd FILL
XFILL_85_DFFSR_243 gnd vdd FILL
XFILL_7_INVX1_4 gnd vdd FILL
XFILL_85_DFFSR_254 gnd vdd FILL
XFILL_85_DFFSR_265 gnd vdd FILL
XFILL_66_7 gnd vdd FILL
XFILL_1_INVX1_160 gnd vdd FILL
XFILL_1_INVX1_171 gnd vdd FILL
XFILL_8_NAND3X1_101 gnd vdd FILL
XFILL_1_INVX1_182 gnd vdd FILL
XFILL_8_NAND3X1_112 gnd vdd FILL
XFILL_1_INVX1_193 gnd vdd FILL
XFILL_8_NAND3X1_123 gnd vdd FILL
XFILL_63_7_2 gnd vdd FILL
XFILL_62_2_1 gnd vdd FILL
XFILL_5_INVX1_170 gnd vdd FILL
XFILL_5_INVX1_181 gnd vdd FILL
XFILL_5_INVX1_192 gnd vdd FILL
XFILL_36_DFFSR_19 gnd vdd FILL
XFILL_76_DFFSR_18 gnd vdd FILL
XFILL_76_DFFSR_29 gnd vdd FILL
XFILL_19_MUX2X1_8 gnd vdd FILL
XFILL_3_NAND2X1_16 gnd vdd FILL
XFILL_3_NAND2X1_27 gnd vdd FILL
XFILL_3_NAND2X1_38 gnd vdd FILL
XFILL_3_NAND2X1_49 gnd vdd FILL
XFILL_0_AND2X2_6 gnd vdd FILL
XFILL_45_DFFSR_17 gnd vdd FILL
XFILL_3_NAND3X1_130 gnd vdd FILL
XFILL_45_DFFSR_28 gnd vdd FILL
XFILL_45_DFFSR_39 gnd vdd FILL
XFILL_13_MUX2X1_180 gnd vdd FILL
XFILL_13_MUX2X1_191 gnd vdd FILL
XFILL_52_DFFSR_210 gnd vdd FILL
XFILL_52_DFFSR_221 gnd vdd FILL
XFILL_52_DFFSR_232 gnd vdd FILL
XFILL_52_DFFSR_243 gnd vdd FILL
XFILL_52_DFFSR_254 gnd vdd FILL
XFILL_85_DFFSR_16 gnd vdd FILL
XFILL_85_DFFSR_27 gnd vdd FILL
XFILL_52_DFFSR_265 gnd vdd FILL
XFILL_12_DFFSR_4 gnd vdd FILL
XFILL_85_DFFSR_38 gnd vdd FILL
XFILL_85_DFFSR_49 gnd vdd FILL
XFILL_29_CLKBUF1_15 gnd vdd FILL
XFILL_14_DFFSR_16 gnd vdd FILL
XFILL_29_CLKBUF1_26 gnd vdd FILL
XFILL_56_DFFSR_220 gnd vdd FILL
XFILL_14_DFFSR_27 gnd vdd FILL
XFILL_14_DFFSR_38 gnd vdd FILL
XFILL_29_CLKBUF1_37 gnd vdd FILL
XFILL_56_DFFSR_231 gnd vdd FILL
XFILL_56_DFFSR_242 gnd vdd FILL
XFILL_14_DFFSR_49 gnd vdd FILL
XFILL_54_7_2 gnd vdd FILL
XFILL_56_DFFSR_253 gnd vdd FILL
XFILL_56_DFFSR_264 gnd vdd FILL
XFILL_56_DFFSR_275 gnd vdd FILL
XFILL_53_2_1 gnd vdd FILL
XFILL_11_CLKBUF1_5 gnd vdd FILL
XFILL_54_DFFSR_15 gnd vdd FILL
XFILL_83_DFFSR_120 gnd vdd FILL
XFILL_7_AOI21X1_16 gnd vdd FILL
XOAI22X1_17 MUX2X1_1/B OAI22X1_4/B INVX1_13/Y OAI22X1_4/D gnd NOR2X1_76/B vdd OAI22X1
XFILL_54_DFFSR_26 gnd vdd FILL
XFILL_83_DFFSR_131 gnd vdd FILL
XFILL_54_DFFSR_37 gnd vdd FILL
XFILL_7_AOI21X1_27 gnd vdd FILL
XOAI22X1_28 INVX1_56/Y OAI22X1_33/B INVX1_61/Y OAI22X1_33/D gnd NOR2X1_89/B vdd OAI22X1
XFILL_83_DFFSR_142 gnd vdd FILL
XFILL_54_DFFSR_48 gnd vdd FILL
XFILL_7_AOI21X1_38 gnd vdd FILL
XFILL_83_DFFSR_153 gnd vdd FILL
XFILL_54_DFFSR_59 gnd vdd FILL
XOAI22X1_39 INVX1_200/Y OAI22X1_49/B INVX1_204/Y OAI22X1_49/D gnd OAI22X1_39/Y vdd
+ OAI22X1
XFILL_7_AOI21X1_49 gnd vdd FILL
XFILL_83_DFFSR_164 gnd vdd FILL
XFILL_83_DFFSR_175 gnd vdd FILL
XFILL_17_OAI22X1_18 gnd vdd FILL
XFILL_15_CLKBUF1_4 gnd vdd FILL
XFILL_3_DFFSR_201 gnd vdd FILL
XFILL_83_DFFSR_186 gnd vdd FILL
XFILL_17_OAI22X1_29 gnd vdd FILL
XFILL_0_NAND3X1_1 gnd vdd FILL
XFILL_83_DFFSR_197 gnd vdd FILL
XFILL_3_DFFSR_212 gnd vdd FILL
XFILL_3_DFFSR_223 gnd vdd FILL
XFILL_87_DFFSR_130 gnd vdd FILL
XFILL_3_DFFSR_234 gnd vdd FILL
XFILL_34_DFFSR_8 gnd vdd FILL
XFILL_3_DFFSR_245 gnd vdd FILL
XFILL_87_DFFSR_141 gnd vdd FILL
XFILL_87_DFFSR_152 gnd vdd FILL
XFILL_23_DFFSR_14 gnd vdd FILL
XFILL_3_DFFSR_256 gnd vdd FILL
XFILL_3_DFFSR_267 gnd vdd FILL
XFILL_23_DFFSR_25 gnd vdd FILL
XFILL_87_DFFSR_163 gnd vdd FILL
XFILL_1_CLKBUF1_19 gnd vdd FILL
XFILL_87_DFFSR_174 gnd vdd FILL
XFILL_19_CLKBUF1_3 gnd vdd FILL
XFILL_7_DFFSR_200 gnd vdd FILL
XFILL_23_DFFSR_36 gnd vdd FILL
XFILL_87_DFFSR_185 gnd vdd FILL
XFILL_23_DFFSR_47 gnd vdd FILL
XFILL_7_DFFSR_211 gnd vdd FILL
XFILL_23_DFFSR_58 gnd vdd FILL
XFILL_87_DFFSR_196 gnd vdd FILL
XFILL_14_BUFX4_90 gnd vdd FILL
XFILL_7_DFFSR_222 gnd vdd FILL
XFILL_23_DFFSR_69 gnd vdd FILL
XFILL_38_DFFSR_209 gnd vdd FILL
XFILL_7_DFFSR_233 gnd vdd FILL
XFILL_7_DFFSR_244 gnd vdd FILL
XFILL_63_DFFSR_13 gnd vdd FILL
XFILL_7_DFFSR_255 gnd vdd FILL
XFILL_63_DFFSR_24 gnd vdd FILL
XFILL_7_DFFSR_266 gnd vdd FILL
XFILL_63_DFFSR_35 gnd vdd FILL
XFILL_63_DFFSR_46 gnd vdd FILL
XFILL_65_DFFSR_109 gnd vdd FILL
XFILL_63_DFFSR_57 gnd vdd FILL
XFILL_63_DFFSR_68 gnd vdd FILL
XFILL_63_DFFSR_79 gnd vdd FILL
XFILL_6_DFFSR_15 gnd vdd FILL
XFILL_6_DFFSR_26 gnd vdd FILL
XFILL_69_DFFSR_108 gnd vdd FILL
XFILL_32_DFFSR_12 gnd vdd FILL
XFILL_6_DFFSR_37 gnd vdd FILL
XFILL_6_DFFSR_48 gnd vdd FILL
XFILL_69_DFFSR_119 gnd vdd FILL
XFILL_32_DFFSR_23 gnd vdd FILL
XFILL_32_DFFSR_34 gnd vdd FILL
XFILL_6_DFFSR_59 gnd vdd FILL
XFILL_32_DFFSR_45 gnd vdd FILL
XFILL_0_AOI22X1_6 gnd vdd FILL
XFILL_32_DFFSR_56 gnd vdd FILL
XFILL_12_OAI21X1_9 gnd vdd FILL
XFILL_7_OAI22X1_13 gnd vdd FILL
XFILL_32_DFFSR_67 gnd vdd FILL
XFILL_7_OAI22X1_24 gnd vdd FILL
XFILL_32_DFFSR_78 gnd vdd FILL
XFILL_7_OAI22X1_35 gnd vdd FILL
XFILL_32_DFFSR_89 gnd vdd FILL
XFILL_7_OAI22X1_46 gnd vdd FILL
XFILL_0_INVX1_205 gnd vdd FILL
XFILL_72_DFFSR_11 gnd vdd FILL
XFILL_45_7_2 gnd vdd FILL
XFILL_72_DFFSR_22 gnd vdd FILL
XFILL_0_INVX1_216 gnd vdd FILL
XFILL_0_INVX1_227 gnd vdd FILL
XFILL_72_DFFSR_33 gnd vdd FILL
XFILL_23_DFFSR_220 gnd vdd FILL
XFILL_72_DFFSR_44 gnd vdd FILL
XFILL_72_DFFSR_55 gnd vdd FILL
XFILL_15_MUX2X1_1 gnd vdd FILL
XFILL_44_2_1 gnd vdd FILL
XFILL_4_AOI22X1_5 gnd vdd FILL
XFILL_23_DFFSR_231 gnd vdd FILL
XFILL_23_DFFSR_242 gnd vdd FILL
XFILL_72_DFFSR_66 gnd vdd FILL
XFILL_72_DFFSR_77 gnd vdd FILL
XFILL_23_DFFSR_253 gnd vdd FILL
XFILL_72_DFFSR_88 gnd vdd FILL
XFILL_23_DFFSR_264 gnd vdd FILL
XFILL_23_DFFSR_275 gnd vdd FILL
XFILL_72_DFFSR_99 gnd vdd FILL
XFILL_4_INVX1_204 gnd vdd FILL
XFILL_4_INVX1_215 gnd vdd FILL
XFILL_50_DFFSR_120 gnd vdd FILL
XFILL_4_INVX1_226 gnd vdd FILL
XFILL_4_NOR2X1_204 gnd vdd FILL
XFILL_50_DFFSR_131 gnd vdd FILL
XFILL_27_DFFSR_230 gnd vdd FILL
XFILL_41_DFFSR_10 gnd vdd FILL
XFILL_8_AOI22X1_4 gnd vdd FILL
XFILL_50_DFFSR_142 gnd vdd FILL
XFILL_27_DFFSR_241 gnd vdd FILL
XFILL_41_DFFSR_21 gnd vdd FILL
XFILL_50_DFFSR_153 gnd vdd FILL
XFILL_27_DFFSR_252 gnd vdd FILL
XFILL_41_DFFSR_32 gnd vdd FILL
XFILL_50_DFFSR_164 gnd vdd FILL
XFILL_41_DFFSR_43 gnd vdd FILL
XFILL_50_DFFSR_175 gnd vdd FILL
XFILL_12_NOR3X1_7 gnd vdd FILL
XFILL_27_DFFSR_263 gnd vdd FILL
XFILL_27_DFFSR_274 gnd vdd FILL
XFILL_0_OAI21X1_15 gnd vdd FILL
XFILL_41_DFFSR_54 gnd vdd FILL
XFILL_50_DFFSR_186 gnd vdd FILL
XFILL_41_DFFSR_65 gnd vdd FILL
XFILL_18_CLKBUF1_11 gnd vdd FILL
XFILL_0_OAI21X1_26 gnd vdd FILL
XFILL_50_DFFSR_197 gnd vdd FILL
XFILL_18_CLKBUF1_22 gnd vdd FILL
XFILL_41_DFFSR_76 gnd vdd FILL
XFILL_0_OAI21X1_37 gnd vdd FILL
XFILL_54_DFFSR_130 gnd vdd FILL
XFILL_18_CLKBUF1_33 gnd vdd FILL
XFILL_41_DFFSR_87 gnd vdd FILL
XFILL_0_OAI21X1_48 gnd vdd FILL
XFILL_41_DFFSR_98 gnd vdd FILL
XFILL_81_DFFSR_20 gnd vdd FILL
XFILL_54_DFFSR_141 gnd vdd FILL
XFILL_54_DFFSR_152 gnd vdd FILL
XFILL_13_AOI21X1_30 gnd vdd FILL
XFILL_54_DFFSR_163 gnd vdd FILL
XFILL_81_DFFSR_31 gnd vdd FILL
XFILL_54_DFFSR_174 gnd vdd FILL
XFILL_81_DFFSR_42 gnd vdd FILL
XFILL_13_AOI21X1_41 gnd vdd FILL
XFILL_81_DFFSR_53 gnd vdd FILL
XFILL_13_AOI21X1_52 gnd vdd FILL
XFILL_10_DFFSR_20 gnd vdd FILL
XFILL_81_DFFSR_64 gnd vdd FILL
XFILL_54_DFFSR_185 gnd vdd FILL
XFILL_81_DFFSR_75 gnd vdd FILL
XFILL_13_AOI21X1_63 gnd vdd FILL
XFILL_54_DFFSR_196 gnd vdd FILL
XFILL_13_AOI21X1_74 gnd vdd FILL
XFILL_10_DFFSR_31 gnd vdd FILL
XFILL_81_DFFSR_86 gnd vdd FILL
XFILL_10_DFFSR_42 gnd vdd FILL
XFILL_10_DFFSR_53 gnd vdd FILL
XFILL_81_DFFSR_97 gnd vdd FILL
XFILL_58_DFFSR_140 gnd vdd FILL
XFILL_10_DFFSR_64 gnd vdd FILL
XFILL_58_DFFSR_151 gnd vdd FILL
XFILL_8_NOR2X1_2 gnd vdd FILL
XFILL_10_DFFSR_75 gnd vdd FILL
XFILL_58_DFFSR_162 gnd vdd FILL
XFILL_10_DFFSR_86 gnd vdd FILL
XFILL_58_DFFSR_173 gnd vdd FILL
XFILL_58_DFFSR_184 gnd vdd FILL
XFILL_1_DFFSR_100 gnd vdd FILL
XFILL_10_DFFSR_97 gnd vdd FILL
XFILL_1_DFFSR_111 gnd vdd FILL
XFILL_32_DFFSR_109 gnd vdd FILL
XFILL_58_DFFSR_195 gnd vdd FILL
XFILL_50_DFFSR_30 gnd vdd FILL
XFILL_1_DFFSR_122 gnd vdd FILL
XFILL_21_NOR3X1_5 gnd vdd FILL
XFILL_1_DFFSR_133 gnd vdd FILL
XFILL_8_2 gnd vdd FILL
XFILL_50_DFFSR_41 gnd vdd FILL
XFILL_1_DFFSR_144 gnd vdd FILL
XFILL_50_DFFSR_52 gnd vdd FILL
XFILL_50_DFFSR_63 gnd vdd FILL
XFILL_1_DFFSR_155 gnd vdd FILL
XFILL_50_DFFSR_74 gnd vdd FILL
XFILL_1_DFFSR_166 gnd vdd FILL
XFILL_50_DFFSR_85 gnd vdd FILL
XFILL_1_DFFSR_177 gnd vdd FILL
XFILL_50_DFFSR_96 gnd vdd FILL
XFILL_1_DFFSR_188 gnd vdd FILL
XFILL_5_DFFSR_110 gnd vdd FILL
XFILL_1_DFFSR_199 gnd vdd FILL
XFILL_36_DFFSR_108 gnd vdd FILL
XFILL_5_DFFSR_121 gnd vdd FILL
XFILL_5_DFFSR_132 gnd vdd FILL
XFILL_36_DFFSR_119 gnd vdd FILL
XFILL_57_3 gnd vdd FILL
XFILL_5_DFFSR_143 gnd vdd FILL
XFILL_5_DFFSR_154 gnd vdd FILL
XFILL_51_DFFSR_2 gnd vdd FILL
XFILL_5_DFFSR_165 gnd vdd FILL
XFILL_36_7_2 gnd vdd FILL
XFILL_5_DFFSR_176 gnd vdd FILL
XFILL_9_NAND3X1_102 gnd vdd FILL
XFILL_9_NAND3X1_113 gnd vdd FILL
XFILL_5_DFFSR_187 gnd vdd FILL
XFILL_5_DFFSR_198 gnd vdd FILL
XFILL_35_2_1 gnd vdd FILL
XFILL_9_NAND3X1_124 gnd vdd FILL
XFILL_9_DFFSR_120 gnd vdd FILL
XFILL_9_DFFSR_131 gnd vdd FILL
XFILL_16_MUX2X1_102 gnd vdd FILL
XFILL_16_MUX2X1_113 gnd vdd FILL
XFILL_9_DFFSR_142 gnd vdd FILL
XFILL_4_NOR3X1_6 gnd vdd FILL
XFILL_13_MUX2X1_40 gnd vdd FILL
XFILL_9_DFFSR_153 gnd vdd FILL
XFILL_16_MUX2X1_124 gnd vdd FILL
XFILL_13_MUX2X1_51 gnd vdd FILL
XFILL_13_MUX2X1_62 gnd vdd FILL
XFILL_9_DFFSR_164 gnd vdd FILL
XFILL_13_MUX2X1_73 gnd vdd FILL
XFILL_9_DFFSR_175 gnd vdd FILL
XFILL_30_NOR3X1_3 gnd vdd FILL
XFILL_16_MUX2X1_135 gnd vdd FILL
XFILL_1_NOR3X1_11 gnd vdd FILL
XFILL_16_MUX2X1_146 gnd vdd FILL
XFILL_13_MUX2X1_84 gnd vdd FILL
XFILL_9_DFFSR_186 gnd vdd FILL
XFILL_1_NOR3X1_22 gnd vdd FILL
XFILL_16_MUX2X1_157 gnd vdd FILL
XFILL_9_DFFSR_197 gnd vdd FILL
XFILL_1_NOR3X1_33 gnd vdd FILL
XFILL_13_MUX2X1_95 gnd vdd FILL
XFILL_16_MUX2X1_168 gnd vdd FILL
XFILL_1_NOR3X1_44 gnd vdd FILL
XFILL_3_AOI21X1_80 gnd vdd FILL
XFILL_16_MUX2X1_179 gnd vdd FILL
XOAI21X1_50 NOR3X1_9/A NOR3X1_9/Y INVX2_2/A gnd OAI21X1_50/Y vdd OAI21X1
XFILL_82_DFFSR_209 gnd vdd FILL
XFILL_17_MUX2X1_50 gnd vdd FILL
XFILL_17_MUX2X1_61 gnd vdd FILL
XFILL_5_NOR3X1_10 gnd vdd FILL
XFILL_17_MUX2X1_72 gnd vdd FILL
XFILL_17_MUX2X1_83 gnd vdd FILL
XFILL_2_DFFSR_30 gnd vdd FILL
XFILL_3_DFFSR_7 gnd vdd FILL
XFILL_2_DFFSR_41 gnd vdd FILL
XFILL_5_NOR3X1_21 gnd vdd FILL
XFILL_16_DFFSR_5 gnd vdd FILL
XFILL_17_MUX2X1_94 gnd vdd FILL
XFILL_5_NOR3X1_32 gnd vdd FILL
XFILL_2_DFFSR_52 gnd vdd FILL
XFILL_5_NOR3X1_43 gnd vdd FILL
XFILL_2_DFFSR_63 gnd vdd FILL
XFILL_73_DFFSR_6 gnd vdd FILL
XFILL_6_NOR2X1_190 gnd vdd FILL
XFILL_2_DFFSR_74 gnd vdd FILL
XFILL_86_DFFSR_208 gnd vdd FILL
XFILL_2_DFFSR_85 gnd vdd FILL
XFILL_21_DFFSR_130 gnd vdd FILL
XFILL_86_DFFSR_219 gnd vdd FILL
XFILL_2_DFFSR_96 gnd vdd FILL
XFILL_21_DFFSR_141 gnd vdd FILL
XFILL_21_DFFSR_152 gnd vdd FILL
XFILL_21_DFFSR_163 gnd vdd FILL
XFILL_21_DFFSR_174 gnd vdd FILL
XFILL_9_NOR3X1_20 gnd vdd FILL
XFILL_9_NOR3X1_31 gnd vdd FILL
XFILL_2_INVX1_103 gnd vdd FILL
XFILL_2_INVX1_114 gnd vdd FILL
XFILL_9_NOR3X1_42 gnd vdd FILL
XFILL_21_DFFSR_185 gnd vdd FILL
XFILL_2_INVX1_125 gnd vdd FILL
XFILL_21_DFFSR_196 gnd vdd FILL
XFILL_2_INVX1_136 gnd vdd FILL
XFILL_2_INVX1_147 gnd vdd FILL
XFILL_25_DFFSR_140 gnd vdd FILL
XFILL_2_INVX1_158 gnd vdd FILL
XFILL_2_INVX1_169 gnd vdd FILL
XFILL_25_DFFSR_151 gnd vdd FILL
XFILL_25_DFFSR_162 gnd vdd FILL
XFILL_25_DFFSR_173 gnd vdd FILL
XFILL_4_NAND3X1_120 gnd vdd FILL
XFILL_25_DFFSR_184 gnd vdd FILL
XFILL_6_INVX1_102 gnd vdd FILL
XFILL_4_NAND3X1_131 gnd vdd FILL
XFILL_23_MUX2X1_170 gnd vdd FILL
XFILL_6_INVX1_113 gnd vdd FILL
XFILL_6_INVX1_124 gnd vdd FILL
XFILL_23_MUX2X1_181 gnd vdd FILL
XFILL_25_DFFSR_195 gnd vdd FILL
XFILL_6_MUX2X1_130 gnd vdd FILL
XFILL_6_INVX1_135 gnd vdd FILL
XFILL_23_MUX2X1_192 gnd vdd FILL
XFILL_6_INVX1_146 gnd vdd FILL
XFILL_6_MUX2X1_141 gnd vdd FILL
XFILL_6_INVX1_157 gnd vdd FILL
XFILL_6_MUX2X1_152 gnd vdd FILL
XFILL_38_DFFSR_9 gnd vdd FILL
XFILL_6_INVX1_168 gnd vdd FILL
XFILL_29_DFFSR_150 gnd vdd FILL
XFILL_29_DFFSR_161 gnd vdd FILL
XFILL_6_MUX2X1_163 gnd vdd FILL
XFILL_6_INVX1_179 gnd vdd FILL
XFILL_29_DFFSR_172 gnd vdd FILL
XFILL_6_MUX2X1_174 gnd vdd FILL
XFILL_6_MUX2X1_185 gnd vdd FILL
XFILL_29_DFFSR_183 gnd vdd FILL
XFILL_29_DFFSR_194 gnd vdd FILL
XFILL_21_NOR3X1_30 gnd vdd FILL
XFILL_21_NOR3X1_41 gnd vdd FILL
XFILL_21_NOR3X1_52 gnd vdd FILL
XFILL_27_7_2 gnd vdd FILL
XFILL_2_7_2 gnd vdd FILL
XFILL_1_2_1 gnd vdd FILL
XFILL_71_DFFSR_230 gnd vdd FILL
XFILL_0_OAI22X1_9 gnd vdd FILL
XFILL_26_2_1 gnd vdd FILL
XFILL_71_DFFSR_241 gnd vdd FILL
XFILL_71_DFFSR_252 gnd vdd FILL
XFILL_71_DFFSR_263 gnd vdd FILL
XFILL_71_DFFSR_274 gnd vdd FILL
XFILL_25_NOR3X1_40 gnd vdd FILL
XFILL_25_NOR3X1_51 gnd vdd FILL
XFILL_4_OAI22X1_8 gnd vdd FILL
XFILL_75_DFFSR_240 gnd vdd FILL
XFILL_10_BUFX4_5 gnd vdd FILL
XFILL_75_DFFSR_251 gnd vdd FILL
XFILL_75_DFFSR_262 gnd vdd FILL
XFILL_30_CLKBUF1_3 gnd vdd FILL
XFILL_75_DFFSR_273 gnd vdd FILL
XFILL_29_NOR3X1_50 gnd vdd FILL
XFILL_10_6_2 gnd vdd FILL
XFILL_8_OAI22X1_7 gnd vdd FILL
XFILL_79_DFFSR_250 gnd vdd FILL
XFILL_79_DFFSR_261 gnd vdd FILL
XFILL_34_CLKBUF1_2 gnd vdd FILL
XFILL_79_DFFSR_272 gnd vdd FILL
XFILL_53_DFFSR_208 gnd vdd FILL
XFILL_9_NAND3X1_11 gnd vdd FILL
XFILL_9_NAND3X1_22 gnd vdd FILL
XFILL_53_DFFSR_219 gnd vdd FILL
XFILL_9_NAND3X1_33 gnd vdd FILL
XFILL_9_NAND3X1_44 gnd vdd FILL
XFILL_9_NAND3X1_55 gnd vdd FILL
XFILL_9_NAND3X1_66 gnd vdd FILL
XFILL_15_BUFX4_13 gnd vdd FILL
XFILL_9_NAND3X1_77 gnd vdd FILL
XFILL_15_BUFX4_24 gnd vdd FILL
XFILL_9_3_1 gnd vdd FILL
XFILL_80_DFFSR_108 gnd vdd FILL
XFILL_15_BUFX4_35 gnd vdd FILL
XFILL_9_NAND3X1_88 gnd vdd FILL
XFILL_57_DFFSR_207 gnd vdd FILL
XFILL_9_NAND3X1_99 gnd vdd FILL
XFILL_15_BUFX4_46 gnd vdd FILL
XFILL_80_DFFSR_119 gnd vdd FILL
XFILL_57_DFFSR_218 gnd vdd FILL
XFILL_15_BUFX4_57 gnd vdd FILL
XFILL_57_DFFSR_229 gnd vdd FILL
XFILL_15_BUFX4_68 gnd vdd FILL
XFILL_15_BUFX4_79 gnd vdd FILL
XFILL_84_DFFSR_107 gnd vdd FILL
XFILL_84_DFFSR_118 gnd vdd FILL
XFILL_84_DFFSR_129 gnd vdd FILL
XFILL_18_7_2 gnd vdd FILL
XFILL_2_NAND2X1_13 gnd vdd FILL
XFILL_2_NAND2X1_24 gnd vdd FILL
XFILL_2_NAND2X1_35 gnd vdd FILL
XFILL_17_2_1 gnd vdd FILL
XFILL_2_NAND2X1_46 gnd vdd FILL
XFILL_2_NAND2X1_57 gnd vdd FILL
XFILL_2_NAND2X1_68 gnd vdd FILL
XFILL_2_NAND2X1_79 gnd vdd FILL
XFILL_13_INVX8_3 gnd vdd FILL
XFILL_60_5_2 gnd vdd FILL
XFILL_5_NAND3X1_9 gnd vdd FILL
XFILL_8_DFFSR_209 gnd vdd FILL
XFILL_42_DFFSR_240 gnd vdd FILL
XFILL_42_DFFSR_251 gnd vdd FILL
XFILL_42_DFFSR_262 gnd vdd FILL
XFILL_42_DFFSR_273 gnd vdd FILL
XFILL_9_NAND3X1_8 gnd vdd FILL
XFILL_28_CLKBUF1_12 gnd vdd FILL
XFILL_28_CLKBUF1_23 gnd vdd FILL
XFILL_55_DFFSR_3 gnd vdd FILL
XFILL_28_CLKBUF1_34 gnd vdd FILL
XFILL_7_BUFX4_12 gnd vdd FILL
XFILL_7_BUFX4_23 gnd vdd FILL
XFILL_46_DFFSR_250 gnd vdd FILL
XFILL_2_AOI22X1_11 gnd vdd FILL
XFILL_7_BUFX4_34 gnd vdd FILL
XFILL_7_BUFX4_45 gnd vdd FILL
XFILL_46_DFFSR_261 gnd vdd FILL
XFILL_46_DFFSR_272 gnd vdd FILL
XFILL_7_BUFX4_56 gnd vdd FILL
XFILL_7_BUFX4_67 gnd vdd FILL
XFILL_20_DFFSR_208 gnd vdd FILL
XFILL_7_BUFX4_78 gnd vdd FILL
XFILL_6_AOI21X1_13 gnd vdd FILL
XFILL_20_DFFSR_219 gnd vdd FILL
XFILL_7_BUFX4_89 gnd vdd FILL
XFILL_6_AOI21X1_24 gnd vdd FILL
XFILL_6_AOI21X1_35 gnd vdd FILL
XFILL_6_AOI21X1_46 gnd vdd FILL
XFILL_73_DFFSR_150 gnd vdd FILL
XFILL_73_DFFSR_161 gnd vdd FILL
XFILL_73_DFFSR_172 gnd vdd FILL
XFILL_16_OAI22X1_15 gnd vdd FILL
XFILL_6_AOI21X1_57 gnd vdd FILL
XFILL_6_AOI21X1_68 gnd vdd FILL
XFILL_73_DFFSR_183 gnd vdd FILL
XFILL_16_OAI22X1_26 gnd vdd FILL
XFILL_6_AOI21X1_79 gnd vdd FILL
XFILL_73_DFFSR_194 gnd vdd FILL
XFILL_16_OAI22X1_37 gnd vdd FILL
XFILL_24_DFFSR_207 gnd vdd FILL
XFILL_9_NOR2X1_101 gnd vdd FILL
XFILL_16_OAI22X1_48 gnd vdd FILL
XFILL_24_DFFSR_218 gnd vdd FILL
XFILL_9_NOR2X1_112 gnd vdd FILL
XFILL_9_NOR2X1_123 gnd vdd FILL
XFILL_24_DFFSR_229 gnd vdd FILL
XFILL_62_1 gnd vdd FILL
XFILL_9_NOR2X1_134 gnd vdd FILL
XFILL_7_DFFSR_8 gnd vdd FILL
XFILL_77_DFFSR_160 gnd vdd FILL
XFILL_9_NOR2X1_145 gnd vdd FILL
XFILL_0_CLKBUF1_16 gnd vdd FILL
XFILL_9_NOR2X1_156 gnd vdd FILL
XFILL_77_DFFSR_171 gnd vdd FILL
XFILL_9_NOR2X1_167 gnd vdd FILL
XFILL_0_CLKBUF1_27 gnd vdd FILL
XFILL_77_DFFSR_182 gnd vdd FILL
XFILL_0_CLKBUF1_38 gnd vdd FILL
XFILL_9_NOR2X1_178 gnd vdd FILL
XFILL_77_DFFSR_193 gnd vdd FILL
XFILL_77_DFFSR_7 gnd vdd FILL
XFILL_51_DFFSR_107 gnd vdd FILL
XFILL_9_NOR2X1_189 gnd vdd FILL
XFILL_28_DFFSR_206 gnd vdd FILL
XFILL_51_DFFSR_118 gnd vdd FILL
XFILL_28_DFFSR_217 gnd vdd FILL
XFILL_15_NAND3X1_80 gnd vdd FILL
XFILL_15_NAND3X1_91 gnd vdd FILL
XFILL_28_DFFSR_228 gnd vdd FILL
XFILL_51_DFFSR_129 gnd vdd FILL
XFILL_51_DFFSR_19 gnd vdd FILL
XFILL_28_DFFSR_239 gnd vdd FILL
XFILL_55_DFFSR_106 gnd vdd FILL
XFILL_55_DFFSR_117 gnd vdd FILL
XFILL_51_5_2 gnd vdd FILL
XFILL_55_DFFSR_128 gnd vdd FILL
XFILL_55_DFFSR_139 gnd vdd FILL
XFILL_50_0_1 gnd vdd FILL
XFILL_20_DFFSR_18 gnd vdd FILL
XFILL_59_DFFSR_105 gnd vdd FILL
XFILL_11_BUFX4_50 gnd vdd FILL
XFILL_20_DFFSR_29 gnd vdd FILL
XFILL_9_MUX2X1_107 gnd vdd FILL
XFILL_9_MUX2X1_118 gnd vdd FILL
XFILL_11_BUFX4_61 gnd vdd FILL
XFILL_59_DFFSR_116 gnd vdd FILL
XFILL_9_MUX2X1_129 gnd vdd FILL
XFILL_59_DFFSR_127 gnd vdd FILL
XFILL_59_DFFSR_138 gnd vdd FILL
XFILL_11_BUFX4_72 gnd vdd FILL
XFILL_11_BUFX4_83 gnd vdd FILL
XFILL_59_DFFSR_149 gnd vdd FILL
XFILL_6_OAI22X1_10 gnd vdd FILL
XFILL_11_BUFX4_94 gnd vdd FILL
XFILL_6_OAI22X1_21 gnd vdd FILL
XFILL_6_OAI22X1_32 gnd vdd FILL
XFILL_6_OAI22X1_43 gnd vdd FILL
XFILL_2_DFFSR_109 gnd vdd FILL
XFILL_60_DFFSR_17 gnd vdd FILL
XDFFSR_20 DFFSR_20/Q DFFSR_88/CLK DFFSR_87/R vdd DFFSR_20/D gnd vdd DFFSR
XFILL_60_DFFSR_28 gnd vdd FILL
XDFFSR_31 DFFSR_31/Q DFFSR_87/CLK DFFSR_87/R vdd DFFSR_31/D gnd vdd DFFSR
XFILL_60_DFFSR_39 gnd vdd FILL
XDFFSR_42 INVX1_18/A DFFSR_56/CLK DFFSR_42/R vdd MUX2X1_5/Y gnd vdd DFFSR
XDFFSR_53 INVX1_11/A DFFSR_81/CLK DFFSR_53/R vdd DFFSR_53/D gnd vdd DFFSR
XDFFSR_64 DFFSR_64/Q DFFSR_64/CLK DFFSR_64/R vdd DFFSR_64/D gnd vdd DFFSR
XDFFSR_75 DFFSR_75/Q DFFSR_78/CLK DFFSR_78/R vdd DFFSR_75/D gnd vdd DFFSR
XFILL_13_DFFSR_250 gnd vdd FILL
XDFFSR_86 DFFSR_86/Q DFFSR_93/CLK DFFSR_93/R vdd DFFSR_86/D gnd vdd DFFSR
XFILL_13_DFFSR_261 gnd vdd FILL
XDFFSR_97 DFFSR_97/Q DFFSR_97/CLK DFFSR_97/R vdd DFFSR_97/D gnd vdd DFFSR
XFILL_6_DFFSR_108 gnd vdd FILL
XFILL_13_DFFSR_272 gnd vdd FILL
XFILL_6_DFFSR_119 gnd vdd FILL
XFILL_10_MUX2X1_17 gnd vdd FILL
XFILL_3_DFFSR_19 gnd vdd FILL
XFILL_10_MUX2X1_28 gnd vdd FILL
XFILL_3_NOR2X1_201 gnd vdd FILL
XFILL_10_MUX2X1_39 gnd vdd FILL
XFILL_1_BUFX4_8 gnd vdd FILL
XFILL_1_AOI21X1_4 gnd vdd FILL
XFILL_40_DFFSR_150 gnd vdd FILL
XFILL_14_BUFX4_6 gnd vdd FILL
XFILL_40_DFFSR_161 gnd vdd FILL
XFILL_17_DFFSR_260 gnd vdd FILL
XFILL_5_INVX1_40 gnd vdd FILL
XFILL_5_NAND3X1_110 gnd vdd FILL
XFILL_59_6_2 gnd vdd FILL
XFILL_40_DFFSR_172 gnd vdd FILL
XFILL_5_NAND3X1_121 gnd vdd FILL
XFILL_17_DFFSR_271 gnd vdd FILL
XFILL_5_NAND3X1_132 gnd vdd FILL
XCLKBUF1_40 BUFX4_4/Y gnd DFFSR_9/CLK vdd CLKBUF1
XFILL_5_INVX1_51 gnd vdd FILL
XFILL_58_1_1 gnd vdd FILL
XFILL_40_DFFSR_183 gnd vdd FILL
XFILL_14_MUX2X1_16 gnd vdd FILL
XFILL_5_INVX1_62 gnd vdd FILL
XFILL_40_DFFSR_194 gnd vdd FILL
XFILL_14_MUX2X1_27 gnd vdd FILL
XFILL_5_INVX1_73 gnd vdd FILL
XFILL_5_INVX1_84 gnd vdd FILL
XFILL_17_CLKBUF1_30 gnd vdd FILL
XFILL_5_INVX1_95 gnd vdd FILL
XFILL_14_MUX2X1_38 gnd vdd FILL
XFILL_17_CLKBUF1_41 gnd vdd FILL
XFILL_5_AOI21X1_3 gnd vdd FILL
XFILL_14_MUX2X1_49 gnd vdd FILL
XFILL_44_DFFSR_160 gnd vdd FILL
XFILL_12_MUX2X1_5 gnd vdd FILL
XFILL_44_DFFSR_171 gnd vdd FILL
XFILL_44_DFFSR_182 gnd vdd FILL
XFILL_18_MUX2X1_15 gnd vdd FILL
XFILL_44_DFFSR_193 gnd vdd FILL
XFILL_12_AOI21X1_60 gnd vdd FILL
XFILL_18_MUX2X1_26 gnd vdd FILL
XFILL_12_AOI21X1_71 gnd vdd FILL
XFILL_18_MUX2X1_37 gnd vdd FILL
XFILL_9_AOI21X1_2 gnd vdd FILL
XFILL_18_MUX2X1_48 gnd vdd FILL
XFILL_18_MUX2X1_59 gnd vdd FILL
XFILL_48_DFFSR_170 gnd vdd FILL
XFILL_3_BUFX4_60 gnd vdd FILL
XFILL_42_5_2 gnd vdd FILL
XFILL_6_NOR3X1_19 gnd vdd FILL
XFILL_3_BUFX4_71 gnd vdd FILL
XFILL_48_DFFSR_181 gnd vdd FILL
XFILL_48_DFFSR_192 gnd vdd FILL
XFILL_3_BUFX4_82 gnd vdd FILL
XFILL_22_DFFSR_106 gnd vdd FILL
XFILL_41_0_1 gnd vdd FILL
XFILL_3_BUFX4_93 gnd vdd FILL
XFILL_22_DFFSR_117 gnd vdd FILL
XFILL_22_DFFSR_128 gnd vdd FILL
XFILL_10_BUFX2_2 gnd vdd FILL
XFILL_22_DFFSR_139 gnd vdd FILL
XFILL_26_DFFSR_105 gnd vdd FILL
XFILL_26_DFFSR_116 gnd vdd FILL
XFILL_21_MUX2X1_3 gnd vdd FILL
XFILL_26_DFFSR_127 gnd vdd FILL
XFILL_26_DFFSR_138 gnd vdd FILL
XFILL_26_DFFSR_149 gnd vdd FILL
XINVX1_103 INVX1_103/A gnd MUX2X1_89/A vdd INVX1
XINVX1_114 DFFSR_90/Q gnd MUX2X1_99/A vdd INVX1
XFILL_5_NOR2X1_6 gnd vdd FILL
XINVX1_125 OAI22X1_7/B gnd INVX1_125/Y vdd INVX1
XINVX1_136 BUFX2_8/A gnd INVX1_136/Y vdd INVX1
XINVX1_147 INVX1_147/A gnd MUX2X1_90/B vdd INVX1
XFILL_29_DFFSR_40 gnd vdd FILL
XFILL_15_MUX2X1_110 gnd vdd FILL
XINVX1_158 INVX1_158/A gnd INVX1_158/Y vdd INVX1
XFILL_15_MUX2X1_121 gnd vdd FILL
XINVX1_169 INVX1_169/A gnd INVX1_169/Y vdd INVX1
XFILL_29_DFFSR_51 gnd vdd FILL
XFILL_15_MUX2X1_132 gnd vdd FILL
XFILL_17_INVX8_4 gnd vdd FILL
XFILL_29_DFFSR_62 gnd vdd FILL
XFILL_29_DFFSR_73 gnd vdd FILL
XFILL_15_MUX2X1_143 gnd vdd FILL
XFILL_29_DFFSR_84 gnd vdd FILL
XFILL_15_MUX2X1_154 gnd vdd FILL
XFILL_15_MUX2X1_165 gnd vdd FILL
XFILL_29_DFFSR_95 gnd vdd FILL
XFILL_22_NOR3X1_17 gnd vdd FILL
XFILL_22_NOR3X1_28 gnd vdd FILL
XFILL_15_MUX2X1_176 gnd vdd FILL
XFILL_15_MUX2X1_187 gnd vdd FILL
XFILL_22_NOR3X1_39 gnd vdd FILL
XFILL_72_DFFSR_206 gnd vdd FILL
XFILL_4_MUX2X1_4 gnd vdd FILL
XFILL_72_DFFSR_217 gnd vdd FILL
XFILL_69_DFFSR_50 gnd vdd FILL
XFILL_72_DFFSR_228 gnd vdd FILL
XFILL_49_1_1 gnd vdd FILL
XFILL_72_DFFSR_239 gnd vdd FILL
XFILL_69_DFFSR_61 gnd vdd FILL
XFILL_69_DFFSR_72 gnd vdd FILL
XFILL_69_DFFSR_83 gnd vdd FILL
XFILL_21_DFFSR_6 gnd vdd FILL
XFILL_26_NOR3X1_16 gnd vdd FILL
XFILL_69_DFFSR_94 gnd vdd FILL
XFILL_26_NOR3X1_27 gnd vdd FILL
XFILL_26_NOR3X1_38 gnd vdd FILL
XFILL_26_NOR3X1_49 gnd vdd FILL
XFILL_76_DFFSR_205 gnd vdd FILL
XFILL_59_DFFSR_4 gnd vdd FILL
XFILL_76_DFFSR_216 gnd vdd FILL
XFILL_76_DFFSR_227 gnd vdd FILL
XFILL_76_DFFSR_238 gnd vdd FILL
XFILL_11_DFFSR_160 gnd vdd FILL
XFILL_76_DFFSR_249 gnd vdd FILL
XFILL_0_CLKBUF1_3 gnd vdd FILL
XFILL_11_DFFSR_171 gnd vdd FILL
XFILL_11_DFFSR_182 gnd vdd FILL
XFILL_38_DFFSR_60 gnd vdd FILL
XFILL_34_5 gnd vdd FILL
XFILL_11_DFFSR_193 gnd vdd FILL
XFILL_38_DFFSR_71 gnd vdd FILL
XFILL_38_DFFSR_82 gnd vdd FILL
XFILL_33_5_2 gnd vdd FILL
XFILL_38_DFFSR_93 gnd vdd FILL
XFILL_27_4 gnd vdd FILL
XFILL_32_0_1 gnd vdd FILL
XFILL_15_DFFSR_170 gnd vdd FILL
XFILL_4_CLKBUF1_2 gnd vdd FILL
XFILL_15_DFFSR_181 gnd vdd FILL
XFILL_15_DFFSR_192 gnd vdd FILL
XFILL_78_DFFSR_70 gnd vdd FILL
XFILL_78_DFFSR_81 gnd vdd FILL
XFILL_78_DFFSR_92 gnd vdd FILL
XFILL_5_MUX2X1_160 gnd vdd FILL
XFILL_8_CLKBUF1_1 gnd vdd FILL
XFILL_5_MUX2X1_171 gnd vdd FILL
XFILL_19_DFFSR_180 gnd vdd FILL
XFILL_5_MUX2X1_182 gnd vdd FILL
XFILL_19_DFFSR_191 gnd vdd FILL
XFILL_5_MUX2X1_193 gnd vdd FILL
XFILL_47_DFFSR_80 gnd vdd FILL
XFILL_47_DFFSR_91 gnd vdd FILL
XFILL_61_DFFSR_260 gnd vdd FILL
XFILL_61_DFFSR_271 gnd vdd FILL
XFILL_87_DFFSR_90 gnd vdd FILL
XFILL_65_DFFSR_270 gnd vdd FILL
XFILL_11_NAND2X1_15 gnd vdd FILL
XFILL_11_NAND2X1_26 gnd vdd FILL
XFILL_16_DFFSR_90 gnd vdd FILL
XFILL_11_NAND2X1_37 gnd vdd FILL
XFILL_11_NAND2X1_48 gnd vdd FILL
XFILL_1_OAI21X1_7 gnd vdd FILL
XFILL_11_NAND2X1_59 gnd vdd FILL
XFILL_43_DFFSR_205 gnd vdd FILL
XFILL_2_NOR2X1_20 gnd vdd FILL
XFILL_2_NOR2X1_31 gnd vdd FILL
XFILL_43_DFFSR_216 gnd vdd FILL
XFILL_2_NOR2X1_42 gnd vdd FILL
XFILL_5_OAI21X1_6 gnd vdd FILL
XFILL_43_DFFSR_227 gnd vdd FILL
XFILL_8_NAND3X1_30 gnd vdd FILL
XFILL_43_DFFSR_238 gnd vdd FILL
XFILL_2_NOR2X1_53 gnd vdd FILL
XFILL_43_DFFSR_249 gnd vdd FILL
XFILL_8_NAND3X1_41 gnd vdd FILL
XFILL_2_NOR2X1_64 gnd vdd FILL
XFILL_8_NAND3X1_52 gnd vdd FILL
XFILL_2_NOR2X1_75 gnd vdd FILL
XFILL_24_5_2 gnd vdd FILL
XFILL_8_NAND3X1_63 gnd vdd FILL
XFILL_8_NAND3X1_74 gnd vdd FILL
XFILL_2_NOR2X1_86 gnd vdd FILL
XFILL_23_0_1 gnd vdd FILL
XFILL_70_DFFSR_105 gnd vdd FILL
XFILL_8_NAND3X1_85 gnd vdd FILL
XFILL_2_NOR2X1_97 gnd vdd FILL
XFILL_47_DFFSR_204 gnd vdd FILL
XFILL_8_NAND3X1_96 gnd vdd FILL
XFILL_70_DFFSR_116 gnd vdd FILL
XFILL_47_DFFSR_215 gnd vdd FILL
XFILL_5_BUFX4_9 gnd vdd FILL
XFILL_9_OAI21X1_5 gnd vdd FILL
XFILL_6_NOR2X1_30 gnd vdd FILL
XFILL_70_DFFSR_127 gnd vdd FILL
XFILL_6_NOR2X1_41 gnd vdd FILL
XFILL_47_DFFSR_226 gnd vdd FILL
XFILL_70_DFFSR_138 gnd vdd FILL
XFILL_6_NOR2X1_52 gnd vdd FILL
XFILL_47_DFFSR_237 gnd vdd FILL
XFILL_70_DFFSR_149 gnd vdd FILL
XFILL_10_OAI22X1_3 gnd vdd FILL
XFILL_47_DFFSR_248 gnd vdd FILL
XFILL_6_NOR2X1_63 gnd vdd FILL
XFILL_47_DFFSR_259 gnd vdd FILL
XFILL_6_NOR2X1_74 gnd vdd FILL
XFILL_6_NOR2X1_85 gnd vdd FILL
XFILL_6_NOR2X1_96 gnd vdd FILL
XFILL_74_DFFSR_104 gnd vdd FILL
XFILL_74_DFFSR_115 gnd vdd FILL
XFILL_74_DFFSR_126 gnd vdd FILL
XFILL_74_DFFSR_137 gnd vdd FILL
XFILL_14_OAI22X1_2 gnd vdd FILL
XFILL_74_DFFSR_148 gnd vdd FILL
XFILL_15_AOI21X1_15 gnd vdd FILL
XFILL_1_NAND2X1_10 gnd vdd FILL
XFILL_15_AOI21X1_26 gnd vdd FILL
XFILL_74_DFFSR_159 gnd vdd FILL
XFILL_15_AOI21X1_37 gnd vdd FILL
XFILL_1_NAND2X1_21 gnd vdd FILL
XFILL_1_NAND2X1_32 gnd vdd FILL
XFILL_15_AOI21X1_48 gnd vdd FILL
XFILL_1_NAND2X1_43 gnd vdd FILL
XFILL_15_AOI21X1_59 gnd vdd FILL
XFILL_78_DFFSR_103 gnd vdd FILL
XFILL_1_NAND2X1_54 gnd vdd FILL
XFILL_78_DFFSR_114 gnd vdd FILL
XFILL_1_NAND2X1_65 gnd vdd FILL
XFILL_12_BUFX4_17 gnd vdd FILL
XFILL_78_DFFSR_125 gnd vdd FILL
XFILL_78_DFFSR_136 gnd vdd FILL
XFILL_12_BUFX4_28 gnd vdd FILL
XFILL_1_NAND2X1_76 gnd vdd FILL
XFILL_1_NAND2X1_87 gnd vdd FILL
XFILL_18_OAI22X1_1 gnd vdd FILL
XFILL_12_BUFX4_39 gnd vdd FILL
XFILL_78_DFFSR_147 gnd vdd FILL
XFILL_78_DFFSR_158 gnd vdd FILL
XFILL_78_DFFSR_169 gnd vdd FILL
XFILL_1_BUFX2_5 gnd vdd FILL
XFILL_7_6_2 gnd vdd FILL
XFILL_6_1_1 gnd vdd FILL
XFILL_6_NAND3X1_100 gnd vdd FILL
XFILL_6_NAND3X1_111 gnd vdd FILL
XFILL_6_NAND3X1_122 gnd vdd FILL
XFILL_32_DFFSR_270 gnd vdd FILL
XFILL_2_NAND2X1_8 gnd vdd FILL
XFILL_27_CLKBUF1_20 gnd vdd FILL
XFILL_60_DFFSR_4 gnd vdd FILL
XFILL_27_CLKBUF1_31 gnd vdd FILL
XFILL_27_CLKBUF1_42 gnd vdd FILL
XFILL_6_INVX1_18 gnd vdd FILL
XFILL_6_NAND2X1_7 gnd vdd FILL
XFILL_10_DFFSR_205 gnd vdd FILL
XFILL_6_INVX1_29 gnd vdd FILL
XFILL_18_MUX2X1_109 gnd vdd FILL
XFILL_5_AOI21X1_10 gnd vdd FILL
XFILL_10_DFFSR_216 gnd vdd FILL
XFILL_15_5_2 gnd vdd FILL
XFILL_5_AOI21X1_21 gnd vdd FILL
XFILL_10_DFFSR_227 gnd vdd FILL
XFILL_2_MUX2X1_60 gnd vdd FILL
XFILL_2_MUX2X1_71 gnd vdd FILL
XFILL_5_AOI21X1_32 gnd vdd FILL
XFILL_10_DFFSR_238 gnd vdd FILL
XFILL_5_AOI21X1_43 gnd vdd FILL
XFILL_2_MUX2X1_82 gnd vdd FILL
XFILL_14_0_1 gnd vdd FILL
XFILL_2_MUX2X1_93 gnd vdd FILL
XFILL_5_AOI21X1_54 gnd vdd FILL
XFILL_10_DFFSR_249 gnd vdd FILL
XFILL_15_OAI22X1_12 gnd vdd FILL
XFILL_63_DFFSR_180 gnd vdd FILL
XFILL_15_OAI22X1_23 gnd vdd FILL
XFILL_5_AOI21X1_65 gnd vdd FILL
XFILL_15_OAI22X1_34 gnd vdd FILL
XFILL_5_AOI21X1_76 gnd vdd FILL
XFILL_63_DFFSR_191 gnd vdd FILL
XFILL_14_DFFSR_204 gnd vdd FILL
XFILL_11_NAND3X1_4 gnd vdd FILL
XFILL_15_OAI22X1_45 gnd vdd FILL
XFILL_14_DFFSR_215 gnd vdd FILL
XFILL_14_DFFSR_226 gnd vdd FILL
XFILL_8_NOR2X1_120 gnd vdd FILL
XFILL_14_DFFSR_237 gnd vdd FILL
XFILL_6_MUX2X1_70 gnd vdd FILL
XFILL_8_NOR2X1_131 gnd vdd FILL
XFILL_6_MUX2X1_81 gnd vdd FILL
XFILL_14_DFFSR_248 gnd vdd FILL
XFILL_8_NOR2X1_142 gnd vdd FILL
XFILL_6_MUX2X1_92 gnd vdd FILL
XFILL_25_DFFSR_7 gnd vdd FILL
XDFFSR_109 INVX1_190/A DFFSR_73/CLK DFFSR_73/R vdd DFFSR_109/D gnd vdd DFFSR
XFILL_4_BUFX4_16 gnd vdd FILL
XFILL_8_NOR2X1_153 gnd vdd FILL
XFILL_14_DFFSR_259 gnd vdd FILL
XFILL_8_NOR2X1_164 gnd vdd FILL
XFILL_4_BUFX4_27 gnd vdd FILL
XFILL_67_DFFSR_190 gnd vdd FILL
XFILL_82_DFFSR_8 gnd vdd FILL
XFILL_8_NOR2X1_175 gnd vdd FILL
XFILL_41_DFFSR_104 gnd vdd FILL
XFILL_18_DFFSR_203 gnd vdd FILL
XFILL_8_NOR2X1_186 gnd vdd FILL
XFILL_4_BUFX4_38 gnd vdd FILL
XFILL_15_NAND3X1_3 gnd vdd FILL
XFILL_8_NOR2X1_197 gnd vdd FILL
XFILL_41_DFFSR_115 gnd vdd FILL
XFILL_4_BUFX4_49 gnd vdd FILL
XFILL_41_DFFSR_126 gnd vdd FILL
XFILL_18_DFFSR_214 gnd vdd FILL
XFILL_18_DFFSR_225 gnd vdd FILL
XFILL_1_INVX2_5 gnd vdd FILL
XFILL_41_DFFSR_137 gnd vdd FILL
XFILL_18_DFFSR_236 gnd vdd FILL
XFILL_41_DFFSR_148 gnd vdd FILL
XFILL_18_DFFSR_247 gnd vdd FILL
XFILL_18_DFFSR_258 gnd vdd FILL
XFILL_41_DFFSR_159 gnd vdd FILL
XFILL_18_DFFSR_269 gnd vdd FILL
XFILL_45_DFFSR_103 gnd vdd FILL
XFILL_45_DFFSR_114 gnd vdd FILL
XFILL_45_DFFSR_125 gnd vdd FILL
XFILL_45_DFFSR_136 gnd vdd FILL
XFILL_45_DFFSR_147 gnd vdd FILL
XFILL_45_DFFSR_158 gnd vdd FILL
XFILL_45_DFFSR_169 gnd vdd FILL
XFILL_8_MUX2X1_104 gnd vdd FILL
XFILL_49_DFFSR_102 gnd vdd FILL
XFILL_8_MUX2X1_115 gnd vdd FILL
XFILL_49_DFFSR_113 gnd vdd FILL
XFILL_49_DFFSR_124 gnd vdd FILL
XFILL_8_MUX2X1_126 gnd vdd FILL
XFILL_49_DFFSR_135 gnd vdd FILL
XFILL_8_MUX2X1_137 gnd vdd FILL
XFILL_49_DFFSR_146 gnd vdd FILL
XFILL_8_MUX2X1_148 gnd vdd FILL
XFILL_11_AND2X2_4 gnd vdd FILL
XFILL_8_MUX2X1_159 gnd vdd FILL
XFILL_49_DFFSR_157 gnd vdd FILL
XFILL_11_AOI22X1_9 gnd vdd FILL
XFILL_49_DFFSR_168 gnd vdd FILL
XFILL_65_4_2 gnd vdd FILL
XFILL_49_DFFSR_179 gnd vdd FILL
XFILL_22_MUX2X1_90 gnd vdd FILL
XFILL_5_OAI22X1_40 gnd vdd FILL
XFILL_5_OAI22X1_51 gnd vdd FILL
XFILL_9_OAI21X1_20 gnd vdd FILL
XFILL_9_OAI21X1_31 gnd vdd FILL
XFILL_9_OAI21X1_42 gnd vdd FILL
XFILL_15_AOI22X1_8 gnd vdd FILL
XFILL_32_2 gnd vdd FILL
XFILL_25_1 gnd vdd FILL
XFILL_19_AOI22X1_7 gnd vdd FILL
XFILL_30_DFFSR_180 gnd vdd FILL
XFILL_39_DFFSR_16 gnd vdd FILL
XFILL_30_DFFSR_191 gnd vdd FILL
XFILL_39_DFFSR_27 gnd vdd FILL
XFILL_39_DFFSR_38 gnd vdd FILL
XFILL_39_DFFSR_49 gnd vdd FILL
XFILL_34_DFFSR_190 gnd vdd FILL
XFILL_79_DFFSR_15 gnd vdd FILL
XFILL_79_DFFSR_26 gnd vdd FILL
XFILL_79_DFFSR_37 gnd vdd FILL
XFILL_79_DFFSR_48 gnd vdd FILL
XFILL_79_DFFSR_59 gnd vdd FILL
XFILL_2_INVX1_11 gnd vdd FILL
XFILL_2_INVX1_22 gnd vdd FILL
XFILL_2_INVX1_33 gnd vdd FILL
XFILL_12_DFFSR_103 gnd vdd FILL
XFILL_2_INVX1_44 gnd vdd FILL
XFILL_12_DFFSR_114 gnd vdd FILL
XFILL_3_AND2X2_3 gnd vdd FILL
XFILL_2_INVX1_55 gnd vdd FILL
XFILL_12_DFFSR_125 gnd vdd FILL
XFILL_2_INVX1_66 gnd vdd FILL
XFILL_12_DFFSR_136 gnd vdd FILL
XFILL_2_INVX1_77 gnd vdd FILL
XFILL_48_DFFSR_14 gnd vdd FILL
XFILL_2_INVX1_88 gnd vdd FILL
XFILL_12_DFFSR_147 gnd vdd FILL
XFILL_12_DFFSR_158 gnd vdd FILL
XFILL_48_DFFSR_25 gnd vdd FILL
XFILL_2_INVX1_99 gnd vdd FILL
XFILL_48_DFFSR_36 gnd vdd FILL
XFILL_12_DFFSR_169 gnd vdd FILL
XFILL_48_DFFSR_47 gnd vdd FILL
XFILL_48_DFFSR_58 gnd vdd FILL
XFILL_16_DFFSR_102 gnd vdd FILL
XFILL_48_DFFSR_69 gnd vdd FILL
XFILL_16_DFFSR_113 gnd vdd FILL
XFILL_16_DFFSR_124 gnd vdd FILL
XFILL_0_NAND3X1_18 gnd vdd FILL
XFILL_56_4_2 gnd vdd FILL
XFILL_16_DFFSR_135 gnd vdd FILL
XFILL_0_NAND3X1_29 gnd vdd FILL
XFILL_16_DFFSR_146 gnd vdd FILL
XFILL_16_DFFSR_157 gnd vdd FILL
XFILL_0_BUFX4_20 gnd vdd FILL
XFILL_42_DFFSR_1 gnd vdd FILL
XFILL_0_BUFX4_31 gnd vdd FILL
XFILL_16_DFFSR_168 gnd vdd FILL
XFILL_16_DFFSR_179 gnd vdd FILL
XFILL_17_DFFSR_13 gnd vdd FILL
XFILL_0_BUFX4_42 gnd vdd FILL
XFILL_17_DFFSR_24 gnd vdd FILL
XFILL_0_BUFX4_53 gnd vdd FILL
XFILL_0_BUFX4_64 gnd vdd FILL
XFILL_17_DFFSR_35 gnd vdd FILL
XFILL_0_BUFX4_75 gnd vdd FILL
XFILL_17_DFFSR_46 gnd vdd FILL
XFILL_0_BUFX4_86 gnd vdd FILL
XFILL_17_DFFSR_57 gnd vdd FILL
XFILL_0_BUFX4_97 gnd vdd FILL
XFILL_17_DFFSR_68 gnd vdd FILL
XFILL_14_MUX2X1_140 gnd vdd FILL
XFILL_17_DFFSR_79 gnd vdd FILL
XFILL_12_NOR3X1_14 gnd vdd FILL
XFILL_14_MUX2X1_151 gnd vdd FILL
XFILL_14_MUX2X1_162 gnd vdd FILL
XFILL_57_DFFSR_12 gnd vdd FILL
XFILL_5_BUFX2_6 gnd vdd FILL
XFILL_14_MUX2X1_173 gnd vdd FILL
XFILL_57_DFFSR_23 gnd vdd FILL
XFILL_12_NOR3X1_25 gnd vdd FILL
XFILL_12_NOR3X1_36 gnd vdd FILL
XFILL_57_DFFSR_34 gnd vdd FILL
XFILL_14_MUX2X1_184 gnd vdd FILL
XFILL_12_NOR3X1_47 gnd vdd FILL
XFILL_28_NOR3X1_9 gnd vdd FILL
XFILL_62_DFFSR_203 gnd vdd FILL
XFILL_57_DFFSR_45 gnd vdd FILL
XFILL_57_DFFSR_56 gnd vdd FILL
XFILL_62_DFFSR_214 gnd vdd FILL
XFILL_57_DFFSR_67 gnd vdd FILL
XFILL_62_DFFSR_225 gnd vdd FILL
XFILL_57_DFFSR_78 gnd vdd FILL
XFILL_62_DFFSR_236 gnd vdd FILL
XFILL_5_BUFX4_105 gnd vdd FILL
XFILL_57_DFFSR_89 gnd vdd FILL
XFILL_62_DFFSR_247 gnd vdd FILL
XFILL_16_NOR3X1_13 gnd vdd FILL
XFILL_62_DFFSR_258 gnd vdd FILL
XFILL_62_DFFSR_269 gnd vdd FILL
XFILL_16_NOR3X1_24 gnd vdd FILL
XFILL_16_NOR3X1_35 gnd vdd FILL
XFILL_66_DFFSR_202 gnd vdd FILL
XFILL_16_NOR3X1_46 gnd vdd FILL
XFILL_64_DFFSR_5 gnd vdd FILL
XFILL_66_DFFSR_213 gnd vdd FILL
XFILL_26_DFFSR_11 gnd vdd FILL
XFILL_9_BUFX4_104 gnd vdd FILL
XFILL_26_DFFSR_22 gnd vdd FILL
XFILL_66_DFFSR_224 gnd vdd FILL
XFILL_66_DFFSR_235 gnd vdd FILL
XFILL_26_DFFSR_33 gnd vdd FILL
XFILL_66_DFFSR_246 gnd vdd FILL
XFILL_26_DFFSR_44 gnd vdd FILL
XFILL_66_DFFSR_257 gnd vdd FILL
XFILL_26_DFFSR_55 gnd vdd FILL
XFILL_66_DFFSR_268 gnd vdd FILL
XFILL_21_CLKBUF1_9 gnd vdd FILL
XFILL_26_DFFSR_66 gnd vdd FILL
XFILL_26_DFFSR_77 gnd vdd FILL
XFILL_26_DFFSR_88 gnd vdd FILL
XFILL_26_DFFSR_99 gnd vdd FILL
XFILL_66_DFFSR_10 gnd vdd FILL
XFILL_66_DFFSR_21 gnd vdd FILL
XFILL_66_DFFSR_32 gnd vdd FILL
XFILL_66_DFFSR_43 gnd vdd FILL
XFILL_1_MUX2X1_8 gnd vdd FILL
XFILL_66_DFFSR_54 gnd vdd FILL
XFILL_25_CLKBUF1_8 gnd vdd FILL
XFILL_66_DFFSR_65 gnd vdd FILL
XFILL_66_DFFSR_76 gnd vdd FILL
XNAND3X1_20 DFFSR_142/Q BUFX4_90/Y AND2X2_4/A gnd OAI21X1_28/C vdd NAND3X1
XFILL_66_DFFSR_87 gnd vdd FILL
XFILL_3_NOR2X1_18 gnd vdd FILL
XFILL_66_DFFSR_98 gnd vdd FILL
XFILL_3_NOR2X1_29 gnd vdd FILL
XNAND3X1_31 AND2X2_7/A INVX1_57/A OAI21X1_41/A gnd NAND3X1_31/Y vdd NAND3X1
XNAND3X1_42 DFFSR_15/Q BUFX4_8/Y NOR2X1_36/Y gnd NAND3X1_46/C vdd NAND3X1
XFILL_9_DFFSR_12 gnd vdd FILL
XNAND3X1_53 NAND3X1_53/A NAND3X1_53/B AOI22X1_5/Y gnd NOR3X1_8/A vdd NAND3X1
XNAND3X1_64 BUFX4_57/Y AND2X2_1/B NOR2X1_42/Y gnd OAI22X1_8/B vdd NAND3X1
XFILL_7_NAND3X1_101 gnd vdd FILL
XFILL_9_DFFSR_23 gnd vdd FILL
XNAND3X1_75 DFFSR_98/Q BUFX4_102/Y NOR2X1_37/Y gnd OAI21X1_6/C vdd NAND3X1
XFILL_29_DFFSR_8 gnd vdd FILL
XFILL_9_DFFSR_34 gnd vdd FILL
XFILL_9_DFFSR_45 gnd vdd FILL
XFILL_7_NAND3X1_112 gnd vdd FILL
XFILL_29_CLKBUF1_7 gnd vdd FILL
XFILL_86_DFFSR_9 gnd vdd FILL
XFILL_47_4_2 gnd vdd FILL
XNAND3X1_86 NOR2X1_4/A BUFX4_7/Y AND2X2_4/A gnd OAI21X1_9/C vdd NAND3X1
XFILL_4_MUX2X1_190 gnd vdd FILL
XFILL_35_DFFSR_20 gnd vdd FILL
XFILL_7_NAND3X1_123 gnd vdd FILL
XFILL_9_DFFSR_56 gnd vdd FILL
XNAND3X1_97 NOR2X1_74/Y NOR3X1_27/Y NOR3X1_18/Y gnd DFFSR_254/D vdd NAND3X1
XFILL_35_DFFSR_31 gnd vdd FILL
XFILL_9_DFFSR_67 gnd vdd FILL
XFILL_35_DFFSR_42 gnd vdd FILL
XNOR2X1_20 NOR2X1_20/A NOR2X1_7/B gnd NOR2X1_20/Y vdd NOR2X1
XFILL_9_DFFSR_78 gnd vdd FILL
XNOR2X1_31 NOR3X1_9/C NOR2X1_37/B gnd NOR2X1_31/Y vdd NOR2X1
XFILL_35_DFFSR_53 gnd vdd FILL
XFILL_7_NOR2X1_17 gnd vdd FILL
XFILL_9_DFFSR_89 gnd vdd FILL
XNOR2X1_42 NOR3X1_9/A NOR3X1_9/B gnd NOR2X1_42/Y vdd NOR2X1
XFILL_7_NOR2X1_28 gnd vdd FILL
XFILL_35_DFFSR_64 gnd vdd FILL
XNOR2X1_53 OAI22X1_2/Y OAI22X1_3/Y gnd NOR2X1_53/Y vdd NOR2X1
XFILL_7_NOR2X1_39 gnd vdd FILL
XFILL_35_DFFSR_75 gnd vdd FILL
XNOR2X1_64 NOR2X1_64/A NOR2X1_64/B gnd NOR2X1_64/Y vdd NOR2X1
XFILL_35_DFFSR_86 gnd vdd FILL
XNOR2X1_75 NOR2X1_75/A NOR2X1_75/B gnd NOR2X1_75/Y vdd NOR2X1
XFILL_35_DFFSR_97 gnd vdd FILL
XNOR2X1_86 INVX1_70/Y NOR2X1_86/B gnd NOR3X1_32/C vdd NOR2X1
XNOR2X1_97 NOR2X1_97/A NOR2X1_97/B gnd NOR2X1_97/Y vdd NOR2X1
XFILL_75_DFFSR_30 gnd vdd FILL
XFILL_75_DFFSR_41 gnd vdd FILL
XFILL_0_NOR2X1_108 gnd vdd FILL
XFILL_75_DFFSR_52 gnd vdd FILL
XFILL_75_DFFSR_63 gnd vdd FILL
XFILL_0_NOR2X1_119 gnd vdd FILL
XFILL_75_DFFSR_74 gnd vdd FILL
XFILL_75_DFFSR_85 gnd vdd FILL
XFILL_3_INVX1_4 gnd vdd FILL
XFILL_75_DFFSR_96 gnd vdd FILL
XFILL_30_3_2 gnd vdd FILL
XFILL_10_NAND2X1_12 gnd vdd FILL
XFILL_10_NAND2X1_23 gnd vdd FILL
XFILL_10_NAND2X1_34 gnd vdd FILL
XFILL_10_NAND2X1_45 gnd vdd FILL
XFILL_15_NOR3X1_4 gnd vdd FILL
XFILL_10_NAND2X1_56 gnd vdd FILL
XFILL_44_DFFSR_40 gnd vdd FILL
XFILL_10_NAND2X1_67 gnd vdd FILL
XFILL_44_DFFSR_51 gnd vdd FILL
XFILL_10_NAND2X1_78 gnd vdd FILL
XFILL_8_OAI22X1_17 gnd vdd FILL
XFILL_44_DFFSR_62 gnd vdd FILL
XFILL_8_OAI22X1_28 gnd vdd FILL
XFILL_10_NAND2X1_89 gnd vdd FILL
XFILL_44_DFFSR_73 gnd vdd FILL
XFILL_8_OAI22X1_39 gnd vdd FILL
XFILL_44_DFFSR_84 gnd vdd FILL
XFILL_33_DFFSR_202 gnd vdd FILL
XFILL_44_DFFSR_95 gnd vdd FILL
XFILL_33_DFFSR_213 gnd vdd FILL
XFILL_33_DFFSR_224 gnd vdd FILL
XFILL_33_DFFSR_235 gnd vdd FILL
XFILL_33_DFFSR_246 gnd vdd FILL
XFILL_84_DFFSR_50 gnd vdd FILL
XFILL_33_DFFSR_257 gnd vdd FILL
XFILL_84_DFFSR_61 gnd vdd FILL
XFILL_2_DFFSR_270 gnd vdd FILL
XFILL_7_NAND3X1_60 gnd vdd FILL
XFILL_2_NAND3X1_130 gnd vdd FILL
XFILL_84_DFFSR_72 gnd vdd FILL
XFILL_84_DFFSR_83 gnd vdd FILL
XFILL_33_DFFSR_268 gnd vdd FILL
XFILL_7_NAND3X1_71 gnd vdd FILL
XFILL_7_NAND3X1_82 gnd vdd FILL
XFILL_84_DFFSR_94 gnd vdd FILL
XFILL_37_DFFSR_201 gnd vdd FILL
XFILL_60_DFFSR_102 gnd vdd FILL
XFILL_13_DFFSR_50 gnd vdd FILL
XFILL_7_NAND3X1_93 gnd vdd FILL
XFILL_37_DFFSR_212 gnd vdd FILL
XFILL_60_DFFSR_113 gnd vdd FILL
XFILL_13_DFFSR_61 gnd vdd FILL
XFILL_60_DFFSR_124 gnd vdd FILL
XFILL_13_DFFSR_72 gnd vdd FILL
XFILL_13_DFFSR_83 gnd vdd FILL
XFILL_60_DFFSR_135 gnd vdd FILL
XFILL_37_DFFSR_223 gnd vdd FILL
XFILL_37_DFFSR_234 gnd vdd FILL
XFILL_13_DFFSR_94 gnd vdd FILL
XFILL_60_DFFSR_146 gnd vdd FILL
XFILL_37_DFFSR_245 gnd vdd FILL
XFILL_60_DFFSR_157 gnd vdd FILL
XFILL_37_DFFSR_256 gnd vdd FILL
XFILL_37_DFFSR_267 gnd vdd FILL
XFILL_60_DFFSR_168 gnd vdd FILL
XFILL_60_DFFSR_179 gnd vdd FILL
XFILL_24_NOR3X1_2 gnd vdd FILL
XFILL_3_MUX2X1_14 gnd vdd FILL
XNAND2X1_8 INVX2_1/A INVX1_68/A gnd NAND2X1_8/Y vdd NAND2X1
XFILL_10_AOI22X1_10 gnd vdd FILL
XFILL_3_MUX2X1_25 gnd vdd FILL
XFILL_1_OAI21X1_19 gnd vdd FILL
XFILL_64_DFFSR_101 gnd vdd FILL
XFILL_3_MUX2X1_36 gnd vdd FILL
XFILL_53_DFFSR_60 gnd vdd FILL
XFILL_19_CLKBUF1_15 gnd vdd FILL
XFILL_64_DFFSR_112 gnd vdd FILL
XFILL_66_7_0 gnd vdd FILL
XFILL_3_MUX2X1_47 gnd vdd FILL
XFILL_19_CLKBUF1_26 gnd vdd FILL
XFILL_53_DFFSR_71 gnd vdd FILL
XFILL_64_DFFSR_123 gnd vdd FILL
XFILL_53_DFFSR_82 gnd vdd FILL
XFILL_64_DFFSR_134 gnd vdd FILL
XFILL_38_4_2 gnd vdd FILL
XFILL_3_MUX2X1_58 gnd vdd FILL
XFILL_19_CLKBUF1_37 gnd vdd FILL
XFILL_3_MUX2X1_69 gnd vdd FILL
XFILL_53_DFFSR_93 gnd vdd FILL
XFILL_64_DFFSR_145 gnd vdd FILL
XFILL_14_AOI21X1_12 gnd vdd FILL
XFILL_64_DFFSR_156 gnd vdd FILL
XFILL_14_AOI21X1_23 gnd vdd FILL
XFILL_14_AOI21X1_34 gnd vdd FILL
XFILL_64_DFFSR_167 gnd vdd FILL
XFILL_14_AOI21X1_45 gnd vdd FILL
XFILL_64_DFFSR_178 gnd vdd FILL
XFILL_7_MUX2X1_13 gnd vdd FILL
XFILL_68_DFFSR_100 gnd vdd FILL
XFILL_64_DFFSR_189 gnd vdd FILL
XFILL_0_NAND2X1_40 gnd vdd FILL
XFILL_7_MUX2X1_24 gnd vdd FILL
XFILL_0_NAND2X1_51 gnd vdd FILL
XFILL_7_MUX2X1_35 gnd vdd FILL
XNOR2X1_110 INVX1_134/A INVX1_137/Y gnd OAI21X1_41/A vdd NOR2X1
XFILL_14_AOI21X1_56 gnd vdd FILL
XFILL_14_AOI21X1_67 gnd vdd FILL
XFILL_0_NAND2X1_62 gnd vdd FILL
XFILL_68_DFFSR_111 gnd vdd FILL
XMUX2X1_60 BUFX4_65/Y INVX1_73/Y NOR2X1_22/Y gnd MUX2X1_60/Y vdd MUX2X1
XNOR2X1_121 INVX1_57/Y NOR2X1_24/B gnd INVX1_205/A vdd NOR2X1
XFILL_7_MUX2X1_46 gnd vdd FILL
XFILL_14_AOI21X1_78 gnd vdd FILL
XNOR2X1_132 DFFSR_140/Q AOI21X1_7/B gnd AOI21X1_5/C vdd NOR2X1
XFILL_68_DFFSR_122 gnd vdd FILL
XFILL_68_DFFSR_133 gnd vdd FILL
XMUX2X1_71 INVX1_84/Y BUFX4_96/Y MUX2X1_71/S gnd MUX2X1_71/Y vdd MUX2X1
XFILL_0_NAND2X1_73 gnd vdd FILL
XFILL_7_MUX2X1_57 gnd vdd FILL
XFILL_68_DFFSR_144 gnd vdd FILL
XNOR2X1_143 NAND2X1_3/Y INVX1_2/Y gnd AOI21X1_9/B vdd NOR2X1
XFILL_7_MUX2X1_68 gnd vdd FILL
XMUX2X1_82 BUFX4_96/Y INVX1_95/Y NOR2X1_28/B gnd MUX2X1_82/Y vdd MUX2X1
XFILL_0_NAND2X1_84 gnd vdd FILL
XFILL_7_MUX2X1_79 gnd vdd FILL
XMUX2X1_93 OAI22X1_7/C BUFX4_64/Y MUX2X1_95/S gnd MUX2X1_93/Y vdd MUX2X1
XFILL_11_OAI21X1_1 gnd vdd FILL
XNOR2X1_154 NAND2X1_3/Y NOR2X1_35/B gnd NOR2X1_154/Y vdd NOR2X1
XFILL_0_NAND2X1_95 gnd vdd FILL
XFILL_68_DFFSR_155 gnd vdd FILL
XNOR2X1_165 NOR2X1_27/A NAND2X1_3/Y gnd NOR2X1_165/Y vdd NOR2X1
XNOR2X1_176 DFFSR_36/Q MUX2X1_14/S gnd NOR2X1_176/Y vdd NOR2X1
XFILL_22_DFFSR_70 gnd vdd FILL
XFILL_68_DFFSR_166 gnd vdd FILL
XFILL_68_DFFSR_177 gnd vdd FILL
XNOR2X1_187 DFFSR_19/Q NOR2X1_190/B gnd NOR2X1_187/Y vdd NOR2X1
XFILL_22_DFFSR_81 gnd vdd FILL
XFILL_22_DFFSR_92 gnd vdd FILL
XFILL_68_DFFSR_188 gnd vdd FILL
XNOR2X1_198 OR2X2_1/B NOR2X1_7/B gnd NOR2X1_202/B vdd NOR2X1
XFILL_7_NOR3X1_3 gnd vdd FILL
XFILL_68_DFFSR_199 gnd vdd FILL
XFILL_21_3_2 gnd vdd FILL
XFILL_62_DFFSR_80 gnd vdd FILL
XFILL_62_DFFSR_91 gnd vdd FILL
XFILL_46_DFFSR_2 gnd vdd FILL
XMUX2X1_105 NAND3X1_30/C INVX1_140/Y AND2X2_8/B gnd OAI21X1_48/B vdd MUX2X1
XFILL_5_DFFSR_60 gnd vdd FILL
XFILL_9_CLKBUF1_10 gnd vdd FILL
XFILL_9_CLKBUF1_21 gnd vdd FILL
XMUX2X1_116 MUX2X1_2/A INVX1_158/Y NOR2X1_128/Y gnd DFFSR_147/D vdd MUX2X1
XFILL_5_DFFSR_71 gnd vdd FILL
XFILL_5_DFFSR_82 gnd vdd FILL
XMUX2X1_127 INVX1_171/Y BUFX4_66/Y NAND2X1_89/Y gnd DFFSR_127/D vdd MUX2X1
XFILL_23_MUX2X1_11 gnd vdd FILL
XFILL_9_CLKBUF1_32 gnd vdd FILL
XFILL_23_MUX2X1_22 gnd vdd FILL
XFILL_5_DFFSR_93 gnd vdd FILL
XMUX2X1_138 BUFX4_93/Y INVX1_182/Y NOR2X1_139/Y gnd DFFSR_120/D vdd MUX2X1
XMUX2X1_149 MUX2X1_1/A INVX1_193/Y NOR2X1_154/Y gnd DFFSR_95/D vdd MUX2X1
XFILL_23_MUX2X1_33 gnd vdd FILL
XFILL_17_MUX2X1_106 gnd vdd FILL
XFILL_23_MUX2X1_44 gnd vdd FILL
XFILL_17_MUX2X1_117 gnd vdd FILL
XFILL_31_DFFSR_90 gnd vdd FILL
XFILL_23_MUX2X1_55 gnd vdd FILL
XFILL_17_MUX2X1_128 gnd vdd FILL
XFILL_23_MUX2X1_66 gnd vdd FILL
XFILL_4_AOI21X1_40 gnd vdd FILL
XFILL_17_MUX2X1_139 gnd vdd FILL
XFILL_23_MUX2X1_77 gnd vdd FILL
XFILL_4_AOI21X1_51 gnd vdd FILL
XFILL_23_MUX2X1_88 gnd vdd FILL
XFILL_4_AOI21X1_62 gnd vdd FILL
XFILL_9_BUFX2_7 gnd vdd FILL
XFILL_23_MUX2X1_99 gnd vdd FILL
XFILL_14_OAI22X1_20 gnd vdd FILL
XFILL_14_OAI22X1_31 gnd vdd FILL
XFILL_4_AOI21X1_73 gnd vdd FILL
XFILL_14_OAI22X1_42 gnd vdd FILL
XINVX1_12 INVX1_12/A gnd NOR3X1_5/A vdd INVX1
XINVX1_23 INVX1_23/A gnd INVX1_23/Y vdd INVX1
XINVX1_34 DFFSR_3/Q gnd INVX1_34/Y vdd INVX1
XINVX1_45 INVX1_45/A gnd INVX1_45/Y vdd INVX1
XINVX1_56 INVX1_56/A gnd INVX1_56/Y vdd INVX1
XFILL_7_NOR2X1_150 gnd vdd FILL
XFILL_30_DFFSR_8 gnd vdd FILL
XINVX1_67 INVX1_67/A gnd NOR3X1_1/A vdd INVX1
XFILL_57_7_0 gnd vdd FILL
XINVX1_78 INVX1_78/A gnd INVX1_78/Y vdd INVX1
XFILL_7_NOR2X1_161 gnd vdd FILL
XFILL_29_4_2 gnd vdd FILL
XINVX1_89 INVX1_89/A gnd INVX1_89/Y vdd INVX1
XFILL_4_4_2 gnd vdd FILL
XFILL_7_NOR2X1_172 gnd vdd FILL
XFILL_31_DFFSR_101 gnd vdd FILL
XFILL_7_NOR2X1_183 gnd vdd FILL
XFILL_68_DFFSR_6 gnd vdd FILL
XFILL_7_NOR2X1_194 gnd vdd FILL
XFILL_31_DFFSR_112 gnd vdd FILL
XFILL_31_DFFSR_123 gnd vdd FILL
XFILL_31_DFFSR_134 gnd vdd FILL
XFILL_31_DFFSR_145 gnd vdd FILL
XFILL_11_NOR2X1_200 gnd vdd FILL
XFILL_31_DFFSR_156 gnd vdd FILL
XFILL_0_DFFSR_180 gnd vdd FILL
XFILL_31_DFFSR_167 gnd vdd FILL
XFILL_31_DFFSR_178 gnd vdd FILL
XFILL_0_DFFSR_191 gnd vdd FILL
XFILL_31_DFFSR_189 gnd vdd FILL
XFILL_35_DFFSR_100 gnd vdd FILL
XFILL_35_DFFSR_111 gnd vdd FILL
XFILL_35_DFFSR_122 gnd vdd FILL
XFILL_35_DFFSR_133 gnd vdd FILL
XFILL_35_DFFSR_144 gnd vdd FILL
XFILL_35_DFFSR_155 gnd vdd FILL
XFILL_35_DFFSR_166 gnd vdd FILL
XFILL_35_DFFSR_177 gnd vdd FILL
XFILL_4_DFFSR_190 gnd vdd FILL
XFILL_40_6_0 gnd vdd FILL
XFILL_35_DFFSR_188 gnd vdd FILL
XFILL_7_MUX2X1_101 gnd vdd FILL
XFILL_12_3_2 gnd vdd FILL
XFILL_7_MUX2X1_112 gnd vdd FILL
XFILL_35_DFFSR_199 gnd vdd FILL
XFILL_39_DFFSR_110 gnd vdd FILL
XFILL_7_MUX2X1_123 gnd vdd FILL
XFILL_39_DFFSR_121 gnd vdd FILL
XFILL_39_DFFSR_132 gnd vdd FILL
XFILL_7_MUX2X1_134 gnd vdd FILL
XFILL_7_MUX2X1_145 gnd vdd FILL
XFILL_39_DFFSR_143 gnd vdd FILL
XFILL_8_BUFX4_1 gnd vdd FILL
XFILL_39_DFFSR_154 gnd vdd FILL
XFILL_7_MUX2X1_156 gnd vdd FILL
XFILL_7_MUX2X1_167 gnd vdd FILL
XFILL_39_DFFSR_165 gnd vdd FILL
XFILL_7_MUX2X1_178 gnd vdd FILL
XFILL_31_NOR3X1_12 gnd vdd FILL
XFILL_39_DFFSR_176 gnd vdd FILL
XFILL_7_MUX2X1_189 gnd vdd FILL
XFILL_39_DFFSR_187 gnd vdd FILL
XFILL_39_DFFSR_198 gnd vdd FILL
XFILL_31_NOR3X1_23 gnd vdd FILL
XFILL_31_NOR3X1_34 gnd vdd FILL
XFILL_81_DFFSR_201 gnd vdd FILL
XFILL_31_NOR3X1_45 gnd vdd FILL
XFILL_8_OAI21X1_50 gnd vdd FILL
XFILL_81_DFFSR_212 gnd vdd FILL
XFILL_81_DFFSR_223 gnd vdd FILL
XFILL_81_DFFSR_234 gnd vdd FILL
XFILL_81_DFFSR_245 gnd vdd FILL
XFILL_81_DFFSR_256 gnd vdd FILL
XFILL_81_DFFSR_267 gnd vdd FILL
XFILL_85_DFFSR_200 gnd vdd FILL
XFILL_85_DFFSR_211 gnd vdd FILL
XFILL_85_DFFSR_222 gnd vdd FILL
XFILL_7_INVX1_5 gnd vdd FILL
XFILL_12_AOI21X1_7 gnd vdd FILL
XFILL_85_DFFSR_233 gnd vdd FILL
XFILL_85_DFFSR_244 gnd vdd FILL
XFILL_85_DFFSR_255 gnd vdd FILL
XFILL_85_DFFSR_266 gnd vdd FILL
XFILL_66_8 gnd vdd FILL
XFILL_48_7_0 gnd vdd FILL
XFILL_1_INVX1_150 gnd vdd FILL
XFILL_1_INVX1_161 gnd vdd FILL
XFILL_8_NAND3X1_102 gnd vdd FILL
XFILL_1_INVX1_172 gnd vdd FILL
XFILL_1_INVX1_183 gnd vdd FILL
XFILL_8_NAND3X1_113 gnd vdd FILL
XFILL_1_INVX1_194 gnd vdd FILL
XFILL_8_NAND3X1_124 gnd vdd FILL
XFILL_62_2_2 gnd vdd FILL
XFILL_5_INVX1_160 gnd vdd FILL
XFILL_5_INVX1_171 gnd vdd FILL
XFILL_5_INVX1_182 gnd vdd FILL
XFILL_8_INVX4_1 gnd vdd FILL
XFILL_5_INVX1_193 gnd vdd FILL
XFILL_31_6_0 gnd vdd FILL
XFILL_76_DFFSR_19 gnd vdd FILL
XFILL_3_NAND2X1_17 gnd vdd FILL
XFILL_19_MUX2X1_9 gnd vdd FILL
XFILL_3_NAND2X1_28 gnd vdd FILL
XFILL_3_NAND2X1_39 gnd vdd FILL
XFILL_0_AND2X2_7 gnd vdd FILL
XFILL_3_NAND3X1_120 gnd vdd FILL
XFILL_45_DFFSR_18 gnd vdd FILL
XFILL_3_NAND3X1_131 gnd vdd FILL
XFILL_13_MUX2X1_170 gnd vdd FILL
XFILL_45_DFFSR_29 gnd vdd FILL
XFILL_13_MUX2X1_181 gnd vdd FILL
XFILL_52_DFFSR_200 gnd vdd FILL
XFILL_13_MUX2X1_192 gnd vdd FILL
XFILL_52_DFFSR_211 gnd vdd FILL
XFILL_52_DFFSR_222 gnd vdd FILL
XFILL_52_DFFSR_233 gnd vdd FILL
XFILL_52_DFFSR_244 gnd vdd FILL
XFILL_52_DFFSR_255 gnd vdd FILL
XFILL_85_DFFSR_17 gnd vdd FILL
XFILL_39_7_0 gnd vdd FILL
XFILL_85_DFFSR_28 gnd vdd FILL
XFILL_12_DFFSR_5 gnd vdd FILL
XFILL_52_DFFSR_266 gnd vdd FILL
XFILL_85_DFFSR_39 gnd vdd FILL
XFILL_56_DFFSR_210 gnd vdd FILL
XFILL_29_CLKBUF1_16 gnd vdd FILL
XFILL_14_DFFSR_17 gnd vdd FILL
XFILL_14_DFFSR_28 gnd vdd FILL
XFILL_29_CLKBUF1_27 gnd vdd FILL
XFILL_29_CLKBUF1_38 gnd vdd FILL
XFILL_56_DFFSR_221 gnd vdd FILL
XFILL_14_DFFSR_39 gnd vdd FILL
XFILL_56_DFFSR_232 gnd vdd FILL
XFILL_56_DFFSR_243 gnd vdd FILL
XFILL_56_DFFSR_254 gnd vdd FILL
XFILL_56_DFFSR_265 gnd vdd FILL
XFILL_53_2_2 gnd vdd FILL
XFILL_11_CLKBUF1_6 gnd vdd FILL
XFILL_54_DFFSR_16 gnd vdd FILL
XFILL_83_DFFSR_110 gnd vdd FILL
XFILL_54_DFFSR_27 gnd vdd FILL
XFILL_83_DFFSR_121 gnd vdd FILL
XOAI22X1_18 INVX1_4/Y OAI22X1_5/B INVX1_9/Y OAI22X1_5/D gnd NOR2X1_77/B vdd OAI22X1
XFILL_83_DFFSR_132 gnd vdd FILL
XFILL_7_AOI21X1_17 gnd vdd FILL
XFILL_54_DFFSR_38 gnd vdd FILL
XFILL_83_DFFSR_143 gnd vdd FILL
XFILL_7_AOI21X1_28 gnd vdd FILL
XOAI22X1_29 INVX1_48/Y OAI22X1_32/B INVX1_52/Y OAI22X1_32/D gnd NOR2X1_89/A vdd OAI22X1
XFILL_7_AOI21X1_39 gnd vdd FILL
XFILL_54_DFFSR_49 gnd vdd FILL
XFILL_83_DFFSR_154 gnd vdd FILL
XFILL_83_DFFSR_165 gnd vdd FILL
XFILL_22_6_0 gnd vdd FILL
XFILL_17_OAI22X1_19 gnd vdd FILL
XFILL_83_DFFSR_176 gnd vdd FILL
XFILL_15_CLKBUF1_5 gnd vdd FILL
XFILL_3_DFFSR_202 gnd vdd FILL
XFILL_83_DFFSR_187 gnd vdd FILL
XFILL_3_DFFSR_213 gnd vdd FILL
XFILL_83_DFFSR_198 gnd vdd FILL
XFILL_0_NAND3X1_2 gnd vdd FILL
XFILL_87_DFFSR_120 gnd vdd FILL
XFILL_3_DFFSR_224 gnd vdd FILL
XFILL_87_DFFSR_131 gnd vdd FILL
XFILL_3_DFFSR_235 gnd vdd FILL
XFILL_87_DFFSR_142 gnd vdd FILL
XFILL_3_DFFSR_246 gnd vdd FILL
XFILL_34_DFFSR_9 gnd vdd FILL
XFILL_87_DFFSR_153 gnd vdd FILL
XFILL_3_DFFSR_257 gnd vdd FILL
XFILL_23_DFFSR_15 gnd vdd FILL
XFILL_11_BUFX4_100 gnd vdd FILL
XFILL_3_DFFSR_268 gnd vdd FILL
XFILL_23_DFFSR_26 gnd vdd FILL
XFILL_87_DFFSR_164 gnd vdd FILL
XFILL_87_DFFSR_175 gnd vdd FILL
XFILL_23_DFFSR_37 gnd vdd FILL
XFILL_19_CLKBUF1_4 gnd vdd FILL
XFILL_7_DFFSR_201 gnd vdd FILL
XFILL_87_DFFSR_186 gnd vdd FILL
XFILL_23_DFFSR_48 gnd vdd FILL
XFILL_14_BUFX4_80 gnd vdd FILL
XFILL_87_DFFSR_197 gnd vdd FILL
XFILL_7_DFFSR_212 gnd vdd FILL
XFILL_4_NAND3X1_1 gnd vdd FILL
XFILL_14_BUFX4_91 gnd vdd FILL
XFILL_23_DFFSR_59 gnd vdd FILL
XFILL_7_DFFSR_223 gnd vdd FILL
XFILL_7_DFFSR_234 gnd vdd FILL
XFILL_7_DFFSR_245 gnd vdd FILL
XDFFSR_270 NOR2X1_9/A DFFSR_9/CLK DFFSR_5/R vdd DFFSR_270/D gnd vdd DFFSR
XFILL_7_DFFSR_256 gnd vdd FILL
XFILL_7_DFFSR_267 gnd vdd FILL
XFILL_63_DFFSR_14 gnd vdd FILL
XFILL_63_DFFSR_25 gnd vdd FILL
XFILL_63_DFFSR_36 gnd vdd FILL
XFILL_63_DFFSR_47 gnd vdd FILL
XFILL_63_DFFSR_58 gnd vdd FILL
XFILL_63_DFFSR_69 gnd vdd FILL
XFILL_6_DFFSR_16 gnd vdd FILL
XFILL_6_DFFSR_27 gnd vdd FILL
XFILL_32_DFFSR_13 gnd vdd FILL
XFILL_6_DFFSR_38 gnd vdd FILL
XFILL_69_DFFSR_109 gnd vdd FILL
XFILL_6_DFFSR_49 gnd vdd FILL
XFILL_32_DFFSR_24 gnd vdd FILL
XFILL_32_DFFSR_35 gnd vdd FILL
XFILL_32_DFFSR_46 gnd vdd FILL
XFILL_5_7_0 gnd vdd FILL
XFILL_32_DFFSR_57 gnd vdd FILL
XFILL_7_OAI22X1_14 gnd vdd FILL
XFILL_0_AOI22X1_7 gnd vdd FILL
XFILL_32_DFFSR_68 gnd vdd FILL
XFILL_7_OAI22X1_25 gnd vdd FILL
XFILL_32_DFFSR_79 gnd vdd FILL
XFILL_7_OAI22X1_36 gnd vdd FILL
XFILL_7_OAI22X1_47 gnd vdd FILL
XFILL_0_INVX1_206 gnd vdd FILL
XFILL_72_DFFSR_12 gnd vdd FILL
XFILL_72_DFFSR_23 gnd vdd FILL
XFILL_23_DFFSR_210 gnd vdd FILL
XFILL_0_INVX1_217 gnd vdd FILL
XFILL_72_DFFSR_34 gnd vdd FILL
XFILL_0_INVX1_228 gnd vdd FILL
XFILL_4_AOI22X1_6 gnd vdd FILL
XFILL_15_MUX2X1_2 gnd vdd FILL
XFILL_23_DFFSR_221 gnd vdd FILL
XFILL_72_DFFSR_45 gnd vdd FILL
XFILL_72_DFFSR_56 gnd vdd FILL
XFILL_44_2_2 gnd vdd FILL
XFILL_23_DFFSR_232 gnd vdd FILL
XFILL_23_DFFSR_243 gnd vdd FILL
XFILL_72_DFFSR_67 gnd vdd FILL
XFILL_72_DFFSR_78 gnd vdd FILL
XFILL_23_DFFSR_254 gnd vdd FILL
XFILL_23_DFFSR_265 gnd vdd FILL
XFILL_72_DFFSR_89 gnd vdd FILL
XFILL_4_INVX1_205 gnd vdd FILL
XFILL_6_NAND3X1_90 gnd vdd FILL
XFILL_4_INVX1_216 gnd vdd FILL
XFILL_50_DFFSR_110 gnd vdd FILL
XFILL_4_NOR2X1_205 gnd vdd FILL
XFILL_27_DFFSR_220 gnd vdd FILL
XFILL_4_INVX1_227 gnd vdd FILL
XFILL_50_DFFSR_121 gnd vdd FILL
XFILL_50_DFFSR_132 gnd vdd FILL
XFILL_8_AOI22X1_5 gnd vdd FILL
XFILL_13_6_0 gnd vdd FILL
XFILL_50_DFFSR_143 gnd vdd FILL
XFILL_41_DFFSR_11 gnd vdd FILL
XFILL_27_DFFSR_231 gnd vdd FILL
XFILL_27_DFFSR_242 gnd vdd FILL
XFILL_41_DFFSR_22 gnd vdd FILL
XFILL_50_DFFSR_154 gnd vdd FILL
XFILL_27_DFFSR_253 gnd vdd FILL
XFILL_41_DFFSR_33 gnd vdd FILL
XFILL_12_NOR3X1_8 gnd vdd FILL
XFILL_6_BUFX4_90 gnd vdd FILL
XFILL_50_DFFSR_165 gnd vdd FILL
XFILL_27_DFFSR_264 gnd vdd FILL
XFILL_50_DFFSR_176 gnd vdd FILL
XFILL_41_DFFSR_44 gnd vdd FILL
XFILL_27_DFFSR_275 gnd vdd FILL
XFILL_41_DFFSR_55 gnd vdd FILL
XFILL_0_OAI21X1_16 gnd vdd FILL
XFILL_50_DFFSR_187 gnd vdd FILL
XFILL_0_OAI21X1_27 gnd vdd FILL
XFILL_41_DFFSR_66 gnd vdd FILL
XFILL_18_CLKBUF1_12 gnd vdd FILL
XFILL_41_DFFSR_77 gnd vdd FILL
XFILL_50_DFFSR_198 gnd vdd FILL
XFILL_0_OAI21X1_38 gnd vdd FILL
XFILL_54_DFFSR_120 gnd vdd FILL
XFILL_18_CLKBUF1_23 gnd vdd FILL
XFILL_41_DFFSR_88 gnd vdd FILL
XFILL_54_DFFSR_131 gnd vdd FILL
XFILL_18_CLKBUF1_34 gnd vdd FILL
XFILL_0_OAI21X1_49 gnd vdd FILL
XFILL_54_DFFSR_142 gnd vdd FILL
XFILL_41_DFFSR_99 gnd vdd FILL
XFILL_81_DFFSR_10 gnd vdd FILL
XFILL_81_DFFSR_21 gnd vdd FILL
XFILL_13_AOI21X1_20 gnd vdd FILL
XFILL_54_DFFSR_153 gnd vdd FILL
XFILL_81_DFFSR_32 gnd vdd FILL
XFILL_81_DFFSR_43 gnd vdd FILL
XFILL_13_AOI21X1_31 gnd vdd FILL
XFILL_54_DFFSR_164 gnd vdd FILL
XFILL_13_AOI21X1_42 gnd vdd FILL
XFILL_54_DFFSR_175 gnd vdd FILL
XFILL_54_DFFSR_186 gnd vdd FILL
XFILL_10_DFFSR_10 gnd vdd FILL
XFILL_81_DFFSR_54 gnd vdd FILL
XFILL_10_DFFSR_21 gnd vdd FILL
XFILL_54_DFFSR_197 gnd vdd FILL
XFILL_81_DFFSR_65 gnd vdd FILL
XFILL_13_AOI21X1_53 gnd vdd FILL
XFILL_81_DFFSR_76 gnd vdd FILL
XFILL_10_DFFSR_32 gnd vdd FILL
XFILL_13_AOI21X1_64 gnd vdd FILL
XFILL_10_DFFSR_43 gnd vdd FILL
XFILL_81_DFFSR_87 gnd vdd FILL
XFILL_13_AOI21X1_75 gnd vdd FILL
XFILL_58_DFFSR_130 gnd vdd FILL
XFILL_81_DFFSR_98 gnd vdd FILL
XFILL_10_DFFSR_54 gnd vdd FILL
XFILL_58_DFFSR_141 gnd vdd FILL
XFILL_58_DFFSR_152 gnd vdd FILL
XFILL_8_NOR2X1_3 gnd vdd FILL
XFILL_10_DFFSR_65 gnd vdd FILL
XFILL_10_DFFSR_76 gnd vdd FILL
XFILL_10_DFFSR_87 gnd vdd FILL
XFILL_58_DFFSR_163 gnd vdd FILL
XFILL_58_DFFSR_174 gnd vdd FILL
XFILL_10_DFFSR_98 gnd vdd FILL
XFILL_1_DFFSR_101 gnd vdd FILL
XFILL_58_DFFSR_185 gnd vdd FILL
XFILL_50_DFFSR_20 gnd vdd FILL
XFILL_1_DFFSR_112 gnd vdd FILL
XFILL_58_DFFSR_196 gnd vdd FILL
XFILL_50_DFFSR_31 gnd vdd FILL
XFILL_1_DFFSR_123 gnd vdd FILL
XFILL_1_DFFSR_134 gnd vdd FILL
XFILL_21_NOR3X1_6 gnd vdd FILL
XFILL_50_DFFSR_42 gnd vdd FILL
XFILL_1_DFFSR_145 gnd vdd FILL
XFILL_8_3 gnd vdd FILL
XFILL_50_DFFSR_53 gnd vdd FILL
XFILL_1_DFFSR_156 gnd vdd FILL
XFILL_50_DFFSR_64 gnd vdd FILL
XFILL_1_DFFSR_167 gnd vdd FILL
XFILL_50_DFFSR_75 gnd vdd FILL
XFILL_1_DFFSR_178 gnd vdd FILL
XFILL_50_DFFSR_86 gnd vdd FILL
XFILL_5_DFFSR_100 gnd vdd FILL
XFILL_1_DFFSR_189 gnd vdd FILL
XFILL_50_DFFSR_97 gnd vdd FILL
XFILL_7_MUX2X1_1 gnd vdd FILL
XFILL_5_DFFSR_111 gnd vdd FILL
XFILL_36_DFFSR_109 gnd vdd FILL
XFILL_5_DFFSR_122 gnd vdd FILL
XFILL_5_DFFSR_133 gnd vdd FILL
XFILL_57_4 gnd vdd FILL
XFILL_5_DFFSR_144 gnd vdd FILL
XFILL_51_DFFSR_3 gnd vdd FILL
XFILL_5_DFFSR_155 gnd vdd FILL
XFILL_5_DFFSR_166 gnd vdd FILL
XFILL_5_DFFSR_177 gnd vdd FILL
XFILL_9_NAND3X1_103 gnd vdd FILL
XFILL_9_NAND3X1_114 gnd vdd FILL
XFILL_5_DFFSR_188 gnd vdd FILL
XFILL_63_5_0 gnd vdd FILL
XFILL_9_DFFSR_110 gnd vdd FILL
XFILL_5_DFFSR_199 gnd vdd FILL
XFILL_35_2_2 gnd vdd FILL
XFILL_9_NAND3X1_125 gnd vdd FILL
XFILL_9_DFFSR_121 gnd vdd FILL
XFILL_16_MUX2X1_103 gnd vdd FILL
XFILL_9_DFFSR_132 gnd vdd FILL
XFILL_13_MUX2X1_30 gnd vdd FILL
XFILL_8_CLKBUF1_40 gnd vdd FILL
XFILL_9_DFFSR_143 gnd vdd FILL
XFILL_13_MUX2X1_41 gnd vdd FILL
XFILL_9_DFFSR_154 gnd vdd FILL
XFILL_16_MUX2X1_114 gnd vdd FILL
XFILL_13_MUX2X1_52 gnd vdd FILL
XFILL_4_NOR3X1_7 gnd vdd FILL
XFILL_16_MUX2X1_125 gnd vdd FILL
XFILL_9_DFFSR_165 gnd vdd FILL
XFILL_16_MUX2X1_136 gnd vdd FILL
XFILL_13_MUX2X1_63 gnd vdd FILL
XFILL_1_NOR3X1_12 gnd vdd FILL
XFILL_13_MUX2X1_74 gnd vdd FILL
XFILL_9_DFFSR_176 gnd vdd FILL
XFILL_30_NOR3X1_4 gnd vdd FILL
XFILL_16_MUX2X1_147 gnd vdd FILL
XFILL_13_MUX2X1_85 gnd vdd FILL
XFILL_9_DFFSR_187 gnd vdd FILL
XFILL_1_NOR3X1_23 gnd vdd FILL
XFILL_3_AOI21X1_70 gnd vdd FILL
XFILL_13_MUX2X1_96 gnd vdd FILL
XFILL_9_DFFSR_198 gnd vdd FILL
XFILL_16_MUX2X1_158 gnd vdd FILL
XFILL_1_NOR3X1_34 gnd vdd FILL
XFILL_16_MUX2X1_169 gnd vdd FILL
XFILL_3_AOI21X1_81 gnd vdd FILL
XOAI21X1_40 INVX2_4/Y INVX2_5/Y AOI22X1_3/A gnd OAI21X1_40/Y vdd OAI21X1
XFILL_1_NOR3X1_45 gnd vdd FILL
XFILL_13_OAI22X1_50 gnd vdd FILL
XFILL_17_MUX2X1_40 gnd vdd FILL
XFILL_17_MUX2X1_51 gnd vdd FILL
XFILL_17_MUX2X1_62 gnd vdd FILL
XFILL_17_MUX2X1_73 gnd vdd FILL
XFILL_5_NOR3X1_11 gnd vdd FILL
XFILL_3_DFFSR_8 gnd vdd FILL
XFILL_2_DFFSR_20 gnd vdd FILL
XFILL_17_MUX2X1_84 gnd vdd FILL
XFILL_2_DFFSR_31 gnd vdd FILL
XFILL_5_NOR3X1_22 gnd vdd FILL
XFILL_17_MUX2X1_95 gnd vdd FILL
XFILL_16_DFFSR_6 gnd vdd FILL
XFILL_2_DFFSR_42 gnd vdd FILL
XFILL_5_NOR3X1_33 gnd vdd FILL
XFILL_2_DFFSR_53 gnd vdd FILL
XFILL_5_NOR3X1_44 gnd vdd FILL
XFILL_6_NOR2X1_180 gnd vdd FILL
XFILL_2_DFFSR_64 gnd vdd FILL
XFILL_6_NOR2X1_191 gnd vdd FILL
XFILL_73_DFFSR_7 gnd vdd FILL
XFILL_21_DFFSR_120 gnd vdd FILL
XFILL_2_DFFSR_75 gnd vdd FILL
XFILL_86_DFFSR_209 gnd vdd FILL
XFILL_21_DFFSR_131 gnd vdd FILL
XFILL_2_DFFSR_86 gnd vdd FILL
XFILL_21_DFFSR_142 gnd vdd FILL
XFILL_2_DFFSR_97 gnd vdd FILL
XFILL_9_NOR3X1_10 gnd vdd FILL
XFILL_21_DFFSR_153 gnd vdd FILL
XFILL_21_DFFSR_164 gnd vdd FILL
XFILL_9_NOR3X1_21 gnd vdd FILL
XFILL_21_DFFSR_175 gnd vdd FILL
XFILL_9_NOR3X1_32 gnd vdd FILL
XFILL_2_INVX1_104 gnd vdd FILL
XFILL_21_DFFSR_186 gnd vdd FILL
XFILL_2_INVX1_115 gnd vdd FILL
XFILL_21_DFFSR_197 gnd vdd FILL
XFILL_9_NOR3X1_43 gnd vdd FILL
XFILL_2_INVX1_126 gnd vdd FILL
XFILL_2_INVX1_137 gnd vdd FILL
XFILL_25_DFFSR_130 gnd vdd FILL
XFILL_2_INVX1_148 gnd vdd FILL
XFILL_25_DFFSR_141 gnd vdd FILL
XFILL_2_INVX1_159 gnd vdd FILL
XFILL_25_DFFSR_152 gnd vdd FILL
XFILL_4_NAND3X1_110 gnd vdd FILL
XFILL_25_DFFSR_163 gnd vdd FILL
XFILL_25_DFFSR_174 gnd vdd FILL
XFILL_4_NAND3X1_121 gnd vdd FILL
XFILL_23_MUX2X1_160 gnd vdd FILL
XFILL_6_INVX1_103 gnd vdd FILL
XFILL_4_NAND3X1_132 gnd vdd FILL
XFILL_25_DFFSR_185 gnd vdd FILL
XFILL_6_INVX1_114 gnd vdd FILL
XFILL_23_MUX2X1_171 gnd vdd FILL
XFILL_25_DFFSR_196 gnd vdd FILL
XFILL_6_INVX1_125 gnd vdd FILL
XFILL_6_MUX2X1_120 gnd vdd FILL
XFILL_23_MUX2X1_182 gnd vdd FILL
XFILL_6_INVX1_136 gnd vdd FILL
XFILL_23_MUX2X1_193 gnd vdd FILL
XFILL_6_INVX1_147 gnd vdd FILL
XFILL_6_MUX2X1_131 gnd vdd FILL
XFILL_29_DFFSR_140 gnd vdd FILL
XFILL_6_MUX2X1_142 gnd vdd FILL
XFILL_6_MUX2X1_153 gnd vdd FILL
XFILL_29_DFFSR_151 gnd vdd FILL
XFILL_6_INVX1_158 gnd vdd FILL
XFILL_29_DFFSR_162 gnd vdd FILL
XFILL_6_INVX1_169 gnd vdd FILL
XFILL_6_MUX2X1_164 gnd vdd FILL
XFILL_6_MUX2X1_175 gnd vdd FILL
XFILL_29_DFFSR_173 gnd vdd FILL
XFILL_29_DFFSR_184 gnd vdd FILL
XFILL_6_MUX2X1_186 gnd vdd FILL
XFILL_21_NOR3X1_20 gnd vdd FILL
XFILL_29_DFFSR_195 gnd vdd FILL
XFILL_21_NOR3X1_31 gnd vdd FILL
XFILL_21_NOR3X1_42 gnd vdd FILL
XFILL_54_5_0 gnd vdd FILL
XFILL_71_DFFSR_220 gnd vdd FILL
XFILL_26_2_2 gnd vdd FILL
XFILL_1_2_2 gnd vdd FILL
XFILL_71_DFFSR_231 gnd vdd FILL
XFILL_71_DFFSR_242 gnd vdd FILL
XFILL_71_DFFSR_253 gnd vdd FILL
XFILL_71_DFFSR_264 gnd vdd FILL
XFILL_25_NOR3X1_30 gnd vdd FILL
XFILL_71_DFFSR_275 gnd vdd FILL
XFILL_25_NOR3X1_41 gnd vdd FILL
XFILL_25_NOR3X1_52 gnd vdd FILL
XFILL_4_OAI22X1_9 gnd vdd FILL
XFILL_75_DFFSR_230 gnd vdd FILL
XFILL_75_DFFSR_241 gnd vdd FILL
XFILL_10_BUFX4_6 gnd vdd FILL
XFILL_75_DFFSR_252 gnd vdd FILL
XFILL_75_DFFSR_263 gnd vdd FILL
XFILL_75_DFFSR_274 gnd vdd FILL
XFILL_30_CLKBUF1_4 gnd vdd FILL
XFILL_29_NOR3X1_40 gnd vdd FILL
XFILL_29_NOR3X1_51 gnd vdd FILL
XFILL_8_OAI22X1_8 gnd vdd FILL
XFILL_79_DFFSR_240 gnd vdd FILL
XFILL_79_DFFSR_251 gnd vdd FILL
XFILL_79_DFFSR_262 gnd vdd FILL
XFILL_34_CLKBUF1_3 gnd vdd FILL
XFILL_79_DFFSR_273 gnd vdd FILL
XFILL_53_DFFSR_209 gnd vdd FILL
XFILL_9_NAND3X1_12 gnd vdd FILL
XFILL_9_NAND3X1_23 gnd vdd FILL
XFILL_9_NAND3X1_34 gnd vdd FILL
XFILL_9_NAND3X1_45 gnd vdd FILL
XFILL_9_NAND3X1_56 gnd vdd FILL
XFILL_9_NAND3X1_67 gnd vdd FILL
XFILL_15_BUFX4_14 gnd vdd FILL
XFILL_9_NAND3X1_78 gnd vdd FILL
XFILL_9_NAND3X1_89 gnd vdd FILL
XFILL_9_3_2 gnd vdd FILL
XFILL_15_BUFX4_25 gnd vdd FILL
XFILL_80_DFFSR_109 gnd vdd FILL
XFILL_57_DFFSR_208 gnd vdd FILL
XFILL_15_BUFX4_36 gnd vdd FILL
XFILL_57_DFFSR_219 gnd vdd FILL
XFILL_15_BUFX4_47 gnd vdd FILL
XFILL_15_BUFX4_58 gnd vdd FILL
XFILL_15_BUFX4_69 gnd vdd FILL
XFILL_84_DFFSR_108 gnd vdd FILL
XFILL_84_DFFSR_119 gnd vdd FILL
XFILL_2_NAND2X1_14 gnd vdd FILL
XFILL_45_5_0 gnd vdd FILL
XFILL_2_NAND2X1_25 gnd vdd FILL
XFILL_2_NAND2X1_36 gnd vdd FILL
XFILL_17_2_2 gnd vdd FILL
XFILL_2_NAND2X1_47 gnd vdd FILL
XFILL_2_NAND2X1_58 gnd vdd FILL
XFILL_2_NAND2X1_69 gnd vdd FILL
XFILL_13_INVX8_4 gnd vdd FILL
XFILL_42_DFFSR_230 gnd vdd FILL
XFILL_42_DFFSR_241 gnd vdd FILL
XFILL_42_DFFSR_252 gnd vdd FILL
XFILL_42_DFFSR_263 gnd vdd FILL
XFILL_42_DFFSR_274 gnd vdd FILL
XFILL_28_CLKBUF1_13 gnd vdd FILL
XFILL_9_NAND3X1_9 gnd vdd FILL
XFILL_28_CLKBUF1_24 gnd vdd FILL
XFILL_55_DFFSR_4 gnd vdd FILL
XFILL_28_CLKBUF1_35 gnd vdd FILL
XFILL_7_BUFX4_13 gnd vdd FILL
XFILL_7_BUFX4_24 gnd vdd FILL
XFILL_46_DFFSR_240 gnd vdd FILL
XFILL_7_BUFX4_35 gnd vdd FILL
XFILL_46_DFFSR_251 gnd vdd FILL
XFILL_46_DFFSR_262 gnd vdd FILL
XFILL_7_BUFX4_46 gnd vdd FILL
XFILL_46_DFFSR_273 gnd vdd FILL
XFILL_7_BUFX4_57 gnd vdd FILL
XFILL_7_BUFX4_68 gnd vdd FILL
XFILL_20_DFFSR_209 gnd vdd FILL
XFILL_7_BUFX4_79 gnd vdd FILL
XFILL_6_AOI21X1_14 gnd vdd FILL
XFILL_73_DFFSR_140 gnd vdd FILL
XFILL_6_AOI21X1_25 gnd vdd FILL
XFILL_73_DFFSR_151 gnd vdd FILL
XFILL_6_AOI21X1_36 gnd vdd FILL
XFILL_6_AOI21X1_47 gnd vdd FILL
XFILL_73_DFFSR_162 gnd vdd FILL
XFILL_6_AOI21X1_58 gnd vdd FILL
XFILL_6_AOI21X1_69 gnd vdd FILL
XFILL_73_DFFSR_173 gnd vdd FILL
XFILL_16_OAI22X1_16 gnd vdd FILL
XFILL_73_DFFSR_184 gnd vdd FILL
XFILL_16_OAI22X1_27 gnd vdd FILL
XFILL_73_DFFSR_195 gnd vdd FILL
XFILL_16_OAI22X1_38 gnd vdd FILL
XFILL_24_DFFSR_208 gnd vdd FILL
XFILL_9_NOR2X1_102 gnd vdd FILL
XFILL_16_OAI22X1_49 gnd vdd FILL
XFILL_9_NOR2X1_113 gnd vdd FILL
XFILL_24_DFFSR_219 gnd vdd FILL
XFILL_9_NOR2X1_124 gnd vdd FILL
XFILL_62_2 gnd vdd FILL
XFILL_7_DFFSR_9 gnd vdd FILL
XFILL_77_DFFSR_150 gnd vdd FILL
XFILL_9_NOR2X1_135 gnd vdd FILL
XFILL_77_DFFSR_161 gnd vdd FILL
XFILL_9_NOR2X1_146 gnd vdd FILL
XFILL_9_NOR2X1_157 gnd vdd FILL
XFILL_0_CLKBUF1_17 gnd vdd FILL
XFILL_77_DFFSR_172 gnd vdd FILL
XFILL_0_CLKBUF1_28 gnd vdd FILL
XFILL_77_DFFSR_183 gnd vdd FILL
XFILL_9_NOR2X1_168 gnd vdd FILL
XFILL_77_DFFSR_8 gnd vdd FILL
XFILL_9_NOR2X1_179 gnd vdd FILL
XFILL_77_DFFSR_194 gnd vdd FILL
XFILL_0_CLKBUF1_39 gnd vdd FILL
XFILL_28_DFFSR_207 gnd vdd FILL
XFILL_51_DFFSR_108 gnd vdd FILL
XFILL_15_NAND3X1_70 gnd vdd FILL
XFILL_15_NAND3X1_81 gnd vdd FILL
XFILL_51_DFFSR_119 gnd vdd FILL
XFILL_28_DFFSR_218 gnd vdd FILL
XFILL_14_AND2X2_1 gnd vdd FILL
XFILL_15_NAND3X1_92 gnd vdd FILL
XFILL_36_5_0 gnd vdd FILL
XFILL_28_DFFSR_229 gnd vdd FILL
XFILL_55_DFFSR_107 gnd vdd FILL
XFILL_55_DFFSR_118 gnd vdd FILL
XFILL_55_DFFSR_129 gnd vdd FILL
XFILL_50_0_2 gnd vdd FILL
XFILL_11_BUFX4_40 gnd vdd FILL
XFILL_20_DFFSR_19 gnd vdd FILL
XFILL_59_DFFSR_106 gnd vdd FILL
XFILL_9_MUX2X1_108 gnd vdd FILL
XFILL_9_MUX2X1_119 gnd vdd FILL
XFILL_11_BUFX4_51 gnd vdd FILL
XFILL_59_DFFSR_117 gnd vdd FILL
XFILL_11_BUFX4_62 gnd vdd FILL
XFILL_11_BUFX4_73 gnd vdd FILL
XFILL_59_DFFSR_128 gnd vdd FILL
XFILL_11_BUFX4_84 gnd vdd FILL
XFILL_59_DFFSR_139 gnd vdd FILL
XFILL_6_OAI22X1_11 gnd vdd FILL
XFILL_11_BUFX4_95 gnd vdd FILL
XFILL_6_OAI22X1_22 gnd vdd FILL
XFILL_6_OAI22X1_33 gnd vdd FILL
XFILL_6_OAI22X1_44 gnd vdd FILL
XDFFSR_10 INVX1_30/A DFFSR_8/CLK DFFSR_8/R vdd DFFSR_10/D gnd vdd DFFSR
XDFFSR_21 DFFSR_21/Q DFFSR_87/CLK DFFSR_93/R vdd DFFSR_21/D gnd vdd DFFSR
XFILL_60_DFFSR_18 gnd vdd FILL
XFILL_60_DFFSR_29 gnd vdd FILL
XDFFSR_32 INVX1_25/A DFFSR_6/CLK DFFSR_6/R vdd DFFSR_32/D gnd vdd DFFSR
XDFFSR_43 INVX1_19/A CLKBUF1_6/Y DFFSR_48/R vdd MUX2X1_6/Y gnd vdd DFFSR
XDFFSR_54 DFFSR_54/Q DFFSR_81/CLK DFFSR_82/R vdd DFFSR_54/D gnd vdd DFFSR
XDFFSR_65 DFFSR_65/Q DFFSR_73/CLK DFFSR_73/R vdd DFFSR_65/D gnd vdd DFFSR
XDFFSR_76 DFFSR_76/Q DFFSR_76/CLK DFFSR_97/R vdd DFFSR_76/D gnd vdd DFFSR
XFILL_13_DFFSR_240 gnd vdd FILL
XFILL_13_DFFSR_251 gnd vdd FILL
XDFFSR_87 DFFSR_87/Q DFFSR_87/CLK DFFSR_87/R vdd DFFSR_87/D gnd vdd DFFSR
XDFFSR_98 DFFSR_98/Q DFFSR_99/CLK DFFSR_98/R vdd DFFSR_98/D gnd vdd DFFSR
XFILL_13_DFFSR_262 gnd vdd FILL
XFILL_13_DFFSR_273 gnd vdd FILL
XFILL_6_DFFSR_109 gnd vdd FILL
XFILL_10_MUX2X1_18 gnd vdd FILL
XFILL_10_MUX2X1_29 gnd vdd FILL
XFILL_3_NOR2X1_202 gnd vdd FILL
XFILL_1_BUFX4_9 gnd vdd FILL
XFILL_1_AOI21X1_5 gnd vdd FILL
XFILL_40_DFFSR_140 gnd vdd FILL
XFILL_40_DFFSR_151 gnd vdd FILL
XFILL_5_NAND3X1_100 gnd vdd FILL
XFILL_14_BUFX4_7 gnd vdd FILL
XFILL_5_INVX1_30 gnd vdd FILL
XFILL_5_NAND3X1_111 gnd vdd FILL
XFILL_17_DFFSR_250 gnd vdd FILL
XFILL_40_DFFSR_162 gnd vdd FILL
XFILL_17_DFFSR_261 gnd vdd FILL
XFILL_5_INVX1_41 gnd vdd FILL
XCLKBUF1_30 BUFX4_10/Y gnd DFFSR_99/CLK vdd CLKBUF1
XFILL_17_DFFSR_272 gnd vdd FILL
XFILL_40_DFFSR_173 gnd vdd FILL
XFILL_5_INVX1_52 gnd vdd FILL
XFILL_5_NAND3X1_122 gnd vdd FILL
XCLKBUF1_41 BUFX4_9/Y gnd DFFSR_45/CLK vdd CLKBUF1
XFILL_40_DFFSR_184 gnd vdd FILL
XFILL_5_INVX1_63 gnd vdd FILL
XFILL_58_1_2 gnd vdd FILL
XFILL_40_DFFSR_195 gnd vdd FILL
XFILL_14_MUX2X1_17 gnd vdd FILL
XFILL_5_INVX1_74 gnd vdd FILL
XFILL_14_MUX2X1_28 gnd vdd FILL
XFILL_17_CLKBUF1_20 gnd vdd FILL
XFILL_5_INVX1_85 gnd vdd FILL
XFILL_14_MUX2X1_39 gnd vdd FILL
XFILL_5_INVX1_96 gnd vdd FILL
XFILL_17_CLKBUF1_31 gnd vdd FILL
XFILL_5_AOI21X1_4 gnd vdd FILL
XFILL_17_CLKBUF1_42 gnd vdd FILL
XFILL_44_DFFSR_150 gnd vdd FILL
XFILL_44_DFFSR_161 gnd vdd FILL
XFILL_12_MUX2X1_6 gnd vdd FILL
XFILL_44_DFFSR_172 gnd vdd FILL
XFILL_12_AOI21X1_50 gnd vdd FILL
XFILL_44_DFFSR_183 gnd vdd FILL
XFILL_27_5_0 gnd vdd FILL
XFILL_18_MUX2X1_16 gnd vdd FILL
XFILL_2_5_0 gnd vdd FILL
XFILL_44_DFFSR_194 gnd vdd FILL
XFILL_18_MUX2X1_27 gnd vdd FILL
XFILL_12_AOI21X1_61 gnd vdd FILL
XFILL_12_AOI21X1_72 gnd vdd FILL
XFILL_18_MUX2X1_38 gnd vdd FILL
XFILL_9_AOI21X1_3 gnd vdd FILL
XFILL_18_MUX2X1_49 gnd vdd FILL
XFILL_10_AOI22X1_1 gnd vdd FILL
XFILL_48_DFFSR_160 gnd vdd FILL
XFILL_3_BUFX4_50 gnd vdd FILL
XFILL_3_BUFX4_61 gnd vdd FILL
XFILL_48_DFFSR_171 gnd vdd FILL
XFILL_3_BUFX4_72 gnd vdd FILL
XFILL_48_DFFSR_182 gnd vdd FILL
XFILL_3_BUFX4_83 gnd vdd FILL
XFILL_41_0_2 gnd vdd FILL
XFILL_48_DFFSR_193 gnd vdd FILL
XFILL_22_DFFSR_107 gnd vdd FILL
XFILL_3_BUFX4_94 gnd vdd FILL
XFILL_22_DFFSR_118 gnd vdd FILL
XFILL_22_DFFSR_129 gnd vdd FILL
XFILL_10_BUFX2_3 gnd vdd FILL
XFILL_10_4_0 gnd vdd FILL
XFILL_26_DFFSR_106 gnd vdd FILL
XFILL_26_DFFSR_117 gnd vdd FILL
XFILL_21_MUX2X1_4 gnd vdd FILL
XFILL_26_DFFSR_128 gnd vdd FILL
XFILL_26_DFFSR_139 gnd vdd FILL
XINVX1_104 INVX1_104/A gnd MUX2X1_91/A vdd INVX1
XFILL_37_DFFSR_1 gnd vdd FILL
XINVX1_115 DFFSR_13/Q gnd NOR3X1_10/A vdd INVX1
XFILL_5_NOR2X1_7 gnd vdd FILL
XINVX1_126 OAI22X1_8/D gnd INVX1_126/Y vdd INVX1
XINVX1_137 INVX1_137/A gnd INVX1_137/Y vdd INVX1
XFILL_15_MUX2X1_100 gnd vdd FILL
XINVX1_148 INVX1_148/A gnd INVX1_148/Y vdd INVX1
XINVX1_159 INVX1_159/A gnd INVX1_159/Y vdd INVX1
XFILL_29_DFFSR_30 gnd vdd FILL
XFILL_15_MUX2X1_111 gnd vdd FILL
XFILL_29_DFFSR_41 gnd vdd FILL
XFILL_15_MUX2X1_122 gnd vdd FILL
XFILL_29_DFFSR_52 gnd vdd FILL
XFILL_29_DFFSR_63 gnd vdd FILL
XFILL_15_MUX2X1_133 gnd vdd FILL
XFILL_15_MUX2X1_144 gnd vdd FILL
XFILL_15_MUX2X1_155 gnd vdd FILL
XFILL_29_DFFSR_74 gnd vdd FILL
XFILL_22_NOR3X1_18 gnd vdd FILL
XFILL_29_DFFSR_85 gnd vdd FILL
XFILL_29_DFFSR_96 gnd vdd FILL
XFILL_15_MUX2X1_166 gnd vdd FILL
XFILL_22_NOR3X1_29 gnd vdd FILL
XFILL_15_MUX2X1_177 gnd vdd FILL
XFILL_15_MUX2X1_188 gnd vdd FILL
XFILL_72_DFFSR_207 gnd vdd FILL
XFILL_69_DFFSR_40 gnd vdd FILL
XFILL_4_MUX2X1_5 gnd vdd FILL
XFILL_72_DFFSR_218 gnd vdd FILL
XFILL_69_DFFSR_51 gnd vdd FILL
XFILL_49_1_2 gnd vdd FILL
XFILL_69_DFFSR_62 gnd vdd FILL
XFILL_72_DFFSR_229 gnd vdd FILL
XFILL_69_DFFSR_73 gnd vdd FILL
XFILL_69_DFFSR_84 gnd vdd FILL
XFILL_26_NOR3X1_17 gnd vdd FILL
XFILL_21_DFFSR_7 gnd vdd FILL
XFILL_69_DFFSR_95 gnd vdd FILL
XFILL_26_NOR3X1_28 gnd vdd FILL
XFILL_26_NOR3X1_39 gnd vdd FILL
XFILL_76_DFFSR_206 gnd vdd FILL
XFILL_59_DFFSR_5 gnd vdd FILL
XFILL_76_DFFSR_217 gnd vdd FILL
XFILL_18_5_0 gnd vdd FILL
XFILL_11_DFFSR_150 gnd vdd FILL
XFILL_76_DFFSR_228 gnd vdd FILL
XFILL_76_DFFSR_239 gnd vdd FILL
XFILL_11_DFFSR_161 gnd vdd FILL
XFILL_11_DFFSR_172 gnd vdd FILL
XFILL_0_CLKBUF1_4 gnd vdd FILL
XFILL_11_DFFSR_183 gnd vdd FILL
XFILL_38_DFFSR_50 gnd vdd FILL
XFILL_11_DFFSR_194 gnd vdd FILL
XFILL_38_DFFSR_61 gnd vdd FILL
XFILL_38_DFFSR_72 gnd vdd FILL
XFILL_38_DFFSR_83 gnd vdd FILL
XFILL_38_DFFSR_94 gnd vdd FILL
XFILL_60_3_0 gnd vdd FILL
XFILL_27_5 gnd vdd FILL
XFILL_15_DFFSR_160 gnd vdd FILL
XFILL_32_0_2 gnd vdd FILL
XFILL_4_CLKBUF1_3 gnd vdd FILL
XFILL_15_DFFSR_171 gnd vdd FILL
XFILL_15_DFFSR_182 gnd vdd FILL
XFILL_15_DFFSR_193 gnd vdd FILL
XFILL_78_DFFSR_60 gnd vdd FILL
XFILL_78_DFFSR_71 gnd vdd FILL
XFILL_78_DFFSR_82 gnd vdd FILL
XFILL_22_MUX2X1_190 gnd vdd FILL
XFILL_78_DFFSR_93 gnd vdd FILL
XFILL_5_MUX2X1_150 gnd vdd FILL
XFILL_5_MUX2X1_161 gnd vdd FILL
XFILL_19_DFFSR_170 gnd vdd FILL
XFILL_5_MUX2X1_172 gnd vdd FILL
XFILL_5_MUX2X1_183 gnd vdd FILL
XFILL_8_CLKBUF1_2 gnd vdd FILL
XFILL_19_DFFSR_181 gnd vdd FILL
XFILL_5_MUX2X1_194 gnd vdd FILL
XFILL_19_DFFSR_192 gnd vdd FILL
XFILL_18_NOR3X1_1 gnd vdd FILL
XFILL_11_NOR3X1_50 gnd vdd FILL
XFILL_47_DFFSR_70 gnd vdd FILL
XFILL_47_DFFSR_81 gnd vdd FILL
XFILL_47_DFFSR_92 gnd vdd FILL
XFILL_61_DFFSR_250 gnd vdd FILL
XFILL_61_DFFSR_261 gnd vdd FILL
XFILL_61_DFFSR_272 gnd vdd FILL
XFILL_87_DFFSR_80 gnd vdd FILL
XFILL_87_DFFSR_91 gnd vdd FILL
XFILL_65_DFFSR_260 gnd vdd FILL
XFILL_65_DFFSR_271 gnd vdd FILL
XFILL_20_CLKBUF1_1 gnd vdd FILL
XFILL_11_NAND2X1_16 gnd vdd FILL
XFILL_16_DFFSR_80 gnd vdd FILL
XFILL_11_NAND2X1_27 gnd vdd FILL
XFILL_16_DFFSR_91 gnd vdd FILL
XFILL_11_NAND2X1_38 gnd vdd FILL
XFILL_11_NAND2X1_49 gnd vdd FILL
XFILL_1_OAI21X1_8 gnd vdd FILL
XFILL_69_DFFSR_270 gnd vdd FILL
XFILL_2_NOR2X1_10 gnd vdd FILL
XFILL_43_DFFSR_206 gnd vdd FILL
XFILL_56_DFFSR_90 gnd vdd FILL
XFILL_43_DFFSR_217 gnd vdd FILL
XFILL_2_NOR2X1_21 gnd vdd FILL
XFILL_8_NAND3X1_20 gnd vdd FILL
XFILL_5_OAI21X1_7 gnd vdd FILL
XFILL_2_NOR2X1_32 gnd vdd FILL
XFILL_2_NOR2X1_43 gnd vdd FILL
XFILL_43_DFFSR_228 gnd vdd FILL
XFILL_8_NAND3X1_31 gnd vdd FILL
XFILL_2_NOR2X1_54 gnd vdd FILL
XFILL_43_DFFSR_239 gnd vdd FILL
XFILL_8_NAND3X1_42 gnd vdd FILL
XFILL_8_NAND3X1_53 gnd vdd FILL
XFILL_2_NOR2X1_65 gnd vdd FILL
XFILL_2_NOR2X1_76 gnd vdd FILL
XFILL_8_NAND3X1_64 gnd vdd FILL
XFILL_51_3_0 gnd vdd FILL
XFILL_8_NAND3X1_75 gnd vdd FILL
XFILL_2_NOR2X1_87 gnd vdd FILL
XFILL_2_NOR2X1_98 gnd vdd FILL
XFILL_8_NAND3X1_86 gnd vdd FILL
XFILL_23_0_2 gnd vdd FILL
XFILL_70_DFFSR_106 gnd vdd FILL
XFILL_47_DFFSR_205 gnd vdd FILL
XFILL_8_NAND3X1_97 gnd vdd FILL
XFILL_6_NOR2X1_20 gnd vdd FILL
XFILL_47_DFFSR_216 gnd vdd FILL
XFILL_70_DFFSR_117 gnd vdd FILL
XFILL_9_OAI21X1_6 gnd vdd FILL
XFILL_6_NOR2X1_31 gnd vdd FILL
XFILL_47_DFFSR_227 gnd vdd FILL
XFILL_70_DFFSR_128 gnd vdd FILL
XFILL_6_NOR2X1_42 gnd vdd FILL
XFILL_70_DFFSR_139 gnd vdd FILL
XFILL_6_NOR2X1_53 gnd vdd FILL
XFILL_10_OAI22X1_4 gnd vdd FILL
XFILL_47_DFFSR_238 gnd vdd FILL
XFILL_47_DFFSR_249 gnd vdd FILL
XFILL_6_NOR2X1_64 gnd vdd FILL
XFILL_6_NOR2X1_75 gnd vdd FILL
XFILL_6_NOR2X1_86 gnd vdd FILL
XFILL_74_DFFSR_105 gnd vdd FILL
XFILL_6_NOR2X1_97 gnd vdd FILL
XFILL_74_DFFSR_116 gnd vdd FILL
XFILL_74_DFFSR_127 gnd vdd FILL
XFILL_74_DFFSR_138 gnd vdd FILL
XFILL_74_DFFSR_149 gnd vdd FILL
XFILL_14_OAI22X1_3 gnd vdd FILL
XFILL_15_AOI21X1_16 gnd vdd FILL
XFILL_1_NAND2X1_11 gnd vdd FILL
XFILL_15_AOI21X1_27 gnd vdd FILL
XFILL_1_NAND2X1_22 gnd vdd FILL
XFILL_15_AOI21X1_38 gnd vdd FILL
XFILL_15_AOI21X1_49 gnd vdd FILL
XFILL_1_NAND2X1_33 gnd vdd FILL
XFILL_78_DFFSR_104 gnd vdd FILL
XFILL_1_NAND2X1_44 gnd vdd FILL
XFILL_1_NAND2X1_55 gnd vdd FILL
XFILL_78_DFFSR_115 gnd vdd FILL
XFILL_1_NAND2X1_66 gnd vdd FILL
XFILL_12_BUFX4_18 gnd vdd FILL
XFILL_1_NAND2X1_77 gnd vdd FILL
XFILL_78_DFFSR_126 gnd vdd FILL
XFILL_78_DFFSR_137 gnd vdd FILL
XFILL_12_BUFX4_29 gnd vdd FILL
XFILL_18_OAI22X1_2 gnd vdd FILL
XFILL_78_DFFSR_148 gnd vdd FILL
XFILL_1_NAND2X1_88 gnd vdd FILL
XFILL_78_DFFSR_159 gnd vdd FILL
XFILL_8_DFFSR_90 gnd vdd FILL
XFILL_1_BUFX2_6 gnd vdd FILL
XFILL_59_4_0 gnd vdd FILL
XFILL_6_NAND3X1_101 gnd vdd FILL
XFILL_6_1_2 gnd vdd FILL
XFILL_6_NAND3X1_112 gnd vdd FILL
XFILL_32_DFFSR_260 gnd vdd FILL
XFILL_32_DFFSR_271 gnd vdd FILL
XFILL_6_NAND3X1_123 gnd vdd FILL
XFILL_27_CLKBUF1_10 gnd vdd FILL
XFILL_2_NAND2X1_9 gnd vdd FILL
XFILL_60_DFFSR_5 gnd vdd FILL
XFILL_27_CLKBUF1_21 gnd vdd FILL
XFILL_27_CLKBUF1_32 gnd vdd FILL
XFILL_36_DFFSR_270 gnd vdd FILL
XFILL_6_INVX1_19 gnd vdd FILL
XFILL_6_NAND2X1_8 gnd vdd FILL
XFILL_10_DFFSR_206 gnd vdd FILL
XFILL_5_AOI21X1_11 gnd vdd FILL
XFILL_2_MUX2X1_50 gnd vdd FILL
XFILL_10_DFFSR_217 gnd vdd FILL
XFILL_5_AOI21X1_22 gnd vdd FILL
XFILL_2_MUX2X1_61 gnd vdd FILL
XFILL_42_3_0 gnd vdd FILL
XFILL_10_DFFSR_228 gnd vdd FILL
XFILL_5_AOI21X1_33 gnd vdd FILL
XFILL_14_0_2 gnd vdd FILL
XFILL_10_DFFSR_239 gnd vdd FILL
XFILL_2_MUX2X1_72 gnd vdd FILL
XFILL_5_AOI21X1_44 gnd vdd FILL
XFILL_2_MUX2X1_83 gnd vdd FILL
XFILL_2_MUX2X1_94 gnd vdd FILL
XFILL_5_AOI21X1_55 gnd vdd FILL
XFILL_63_DFFSR_170 gnd vdd FILL
XFILL_5_AOI21X1_66 gnd vdd FILL
XFILL_15_OAI22X1_13 gnd vdd FILL
XFILL_5_AOI21X1_77 gnd vdd FILL
XFILL_15_OAI22X1_24 gnd vdd FILL
XFILL_63_DFFSR_181 gnd vdd FILL
XFILL_15_OAI22X1_35 gnd vdd FILL
XFILL_63_DFFSR_192 gnd vdd FILL
XFILL_14_DFFSR_205 gnd vdd FILL
XFILL_15_OAI22X1_46 gnd vdd FILL
XFILL_14_DFFSR_216 gnd vdd FILL
XFILL_8_NOR2X1_110 gnd vdd FILL
XFILL_11_NAND3X1_5 gnd vdd FILL
XFILL_6_MUX2X1_60 gnd vdd FILL
XFILL_6_MUX2X1_71 gnd vdd FILL
XFILL_14_DFFSR_227 gnd vdd FILL
XFILL_8_NOR2X1_121 gnd vdd FILL
XFILL_8_NOR2X1_132 gnd vdd FILL
XFILL_14_DFFSR_238 gnd vdd FILL
XFILL_8_NOR2X1_143 gnd vdd FILL
XFILL_14_DFFSR_249 gnd vdd FILL
XFILL_6_MUX2X1_82 gnd vdd FILL
XFILL_6_MUX2X1_93 gnd vdd FILL
XFILL_25_DFFSR_8 gnd vdd FILL
XFILL_8_NOR2X1_154 gnd vdd FILL
XFILL_4_BUFX4_17 gnd vdd FILL
XFILL_8_NOR2X1_165 gnd vdd FILL
XFILL_82_DFFSR_9 gnd vdd FILL
XFILL_67_DFFSR_180 gnd vdd FILL
XFILL_4_BUFX4_28 gnd vdd FILL
XFILL_8_NOR2X1_176 gnd vdd FILL
XFILL_4_BUFX4_39 gnd vdd FILL
XFILL_67_DFFSR_191 gnd vdd FILL
XFILL_8_NOR2X1_187 gnd vdd FILL
XFILL_41_DFFSR_105 gnd vdd FILL
XFILL_18_DFFSR_204 gnd vdd FILL
XFILL_18_DFFSR_215 gnd vdd FILL
XFILL_8_NOR2X1_198 gnd vdd FILL
XFILL_41_DFFSR_116 gnd vdd FILL
XFILL_15_NAND3X1_4 gnd vdd FILL
XFILL_41_DFFSR_127 gnd vdd FILL
XFILL_18_DFFSR_226 gnd vdd FILL
XFILL_41_DFFSR_138 gnd vdd FILL
XFILL_41_DFFSR_149 gnd vdd FILL
XFILL_18_DFFSR_237 gnd vdd FILL
XFILL_18_DFFSR_248 gnd vdd FILL
XFILL_18_DFFSR_259 gnd vdd FILL
XFILL_1_NAND3X1_130 gnd vdd FILL
XFILL_45_DFFSR_104 gnd vdd FILL
XFILL_45_DFFSR_115 gnd vdd FILL
XFILL_45_DFFSR_126 gnd vdd FILL
XFILL_45_DFFSR_137 gnd vdd FILL
XFILL_45_DFFSR_148 gnd vdd FILL
XFILL_45_DFFSR_159 gnd vdd FILL
XFILL_49_DFFSR_103 gnd vdd FILL
XFILL_8_MUX2X1_105 gnd vdd FILL
XFILL_8_MUX2X1_116 gnd vdd FILL
XFILL_49_DFFSR_114 gnd vdd FILL
XFILL_8_MUX2X1_127 gnd vdd FILL
XFILL_49_DFFSR_125 gnd vdd FILL
XFILL_49_DFFSR_136 gnd vdd FILL
XFILL_8_MUX2X1_138 gnd vdd FILL
XFILL_8_MUX2X1_149 gnd vdd FILL
XFILL_49_DFFSR_147 gnd vdd FILL
XFILL_49_DFFSR_158 gnd vdd FILL
XFILL_11_AND2X2_5 gnd vdd FILL
XFILL_5_OAI22X1_30 gnd vdd FILL
XFILL_49_DFFSR_169 gnd vdd FILL
XFILL_22_MUX2X1_80 gnd vdd FILL
XFILL_22_MUX2X1_91 gnd vdd FILL
XFILL_5_OAI22X1_41 gnd vdd FILL
XFILL_9_OAI21X1_10 gnd vdd FILL
XFILL_9_OAI21X1_21 gnd vdd FILL
XFILL_9_OAI21X1_32 gnd vdd FILL
XFILL_9_OAI21X1_43 gnd vdd FILL
XFILL_15_AOI22X1_9 gnd vdd FILL
XFILL_32_3 gnd vdd FILL
XFILL_33_3_0 gnd vdd FILL
XFILL_25_2 gnd vdd FILL
XFILL_19_AOI22X1_8 gnd vdd FILL
XFILL_18_1 gnd vdd FILL
XFILL_30_DFFSR_170 gnd vdd FILL
XFILL_30_DFFSR_181 gnd vdd FILL
XFILL_39_DFFSR_17 gnd vdd FILL
XFILL_30_DFFSR_192 gnd vdd FILL
XFILL_39_DFFSR_28 gnd vdd FILL
XFILL_39_DFFSR_39 gnd vdd FILL
XFILL_34_DFFSR_180 gnd vdd FILL
XFILL_79_DFFSR_16 gnd vdd FILL
XFILL_34_DFFSR_191 gnd vdd FILL
XFILL_79_DFFSR_27 gnd vdd FILL
XFILL_79_DFFSR_38 gnd vdd FILL
XFILL_11_AOI21X1_80 gnd vdd FILL
XFILL_79_DFFSR_49 gnd vdd FILL
XFILL_2_INVX1_12 gnd vdd FILL
XFILL_2_INVX1_23 gnd vdd FILL
XFILL_2_INVX1_34 gnd vdd FILL
XFILL_12_DFFSR_104 gnd vdd FILL
XFILL_38_DFFSR_190 gnd vdd FILL
XFILL_3_AND2X2_4 gnd vdd FILL
XFILL_2_INVX1_45 gnd vdd FILL
XFILL_2_INVX1_56 gnd vdd FILL
XFILL_12_DFFSR_115 gnd vdd FILL
XFILL_2_INVX1_67 gnd vdd FILL
XFILL_12_DFFSR_126 gnd vdd FILL
XFILL_12_DFFSR_137 gnd vdd FILL
XFILL_12_DFFSR_148 gnd vdd FILL
XFILL_2_INVX1_78 gnd vdd FILL
XFILL_48_DFFSR_15 gnd vdd FILL
XFILL_2_INVX1_89 gnd vdd FILL
XFILL_48_DFFSR_26 gnd vdd FILL
XFILL_48_DFFSR_37 gnd vdd FILL
XFILL_12_DFFSR_159 gnd vdd FILL
XFILL_48_DFFSR_48 gnd vdd FILL
XFILL_80_DFFSR_270 gnd vdd FILL
XFILL_16_DFFSR_103 gnd vdd FILL
XFILL_48_DFFSR_59 gnd vdd FILL
XFILL_16_DFFSR_114 gnd vdd FILL
XFILL_0_NAND3X1_19 gnd vdd FILL
XFILL_16_DFFSR_125 gnd vdd FILL
XFILL_16_DFFSR_136 gnd vdd FILL
XFILL_16_DFFSR_147 gnd vdd FILL
XFILL_0_BUFX4_10 gnd vdd FILL
XFILL_16_DFFSR_158 gnd vdd FILL
XFILL_0_BUFX4_21 gnd vdd FILL
XFILL_42_DFFSR_2 gnd vdd FILL
XFILL_16_DFFSR_169 gnd vdd FILL
XFILL_0_BUFX4_32 gnd vdd FILL
XFILL_0_BUFX4_43 gnd vdd FILL
XFILL_0_BUFX4_54 gnd vdd FILL
XFILL_17_DFFSR_14 gnd vdd FILL
XFILL_17_DFFSR_25 gnd vdd FILL
XFILL_17_DFFSR_36 gnd vdd FILL
XFILL_0_BUFX4_65 gnd vdd FILL
XFILL_0_BUFX4_76 gnd vdd FILL
XFILL_17_DFFSR_47 gnd vdd FILL
XFILL_0_BUFX4_87 gnd vdd FILL
XFILL_17_DFFSR_58 gnd vdd FILL
XFILL_0_BUFX4_98 gnd vdd FILL
XFILL_17_DFFSR_69 gnd vdd FILL
XFILL_14_MUX2X1_130 gnd vdd FILL
XFILL_24_3_0 gnd vdd FILL
XFILL_14_MUX2X1_141 gnd vdd FILL
XFILL_14_MUX2X1_152 gnd vdd FILL
XFILL_14_MUX2X1_163 gnd vdd FILL
XFILL_12_NOR3X1_15 gnd vdd FILL
XFILL_57_DFFSR_13 gnd vdd FILL
XFILL_12_NOR3X1_26 gnd vdd FILL
XFILL_5_BUFX2_7 gnd vdd FILL
XFILL_57_DFFSR_24 gnd vdd FILL
XFILL_14_MUX2X1_174 gnd vdd FILL
XFILL_57_DFFSR_35 gnd vdd FILL
XFILL_14_MUX2X1_185 gnd vdd FILL
XFILL_12_NOR3X1_37 gnd vdd FILL
XFILL_57_DFFSR_46 gnd vdd FILL
XFILL_12_NOR3X1_48 gnd vdd FILL
XFILL_62_DFFSR_204 gnd vdd FILL
XFILL_62_DFFSR_215 gnd vdd FILL
XFILL_57_DFFSR_57 gnd vdd FILL
XFILL_62_DFFSR_226 gnd vdd FILL
XFILL_57_DFFSR_68 gnd vdd FILL
XFILL_62_DFFSR_237 gnd vdd FILL
XFILL_57_DFFSR_79 gnd vdd FILL
XFILL_62_DFFSR_248 gnd vdd FILL
XFILL_16_NOR3X1_14 gnd vdd FILL
XFILL_62_DFFSR_259 gnd vdd FILL
XFILL_16_NOR3X1_25 gnd vdd FILL
XFILL_16_NOR3X1_36 gnd vdd FILL
XFILL_16_NOR3X1_47 gnd vdd FILL
XFILL_66_DFFSR_203 gnd vdd FILL
XFILL_26_DFFSR_12 gnd vdd FILL
XFILL_64_DFFSR_6 gnd vdd FILL
XFILL_66_DFFSR_214 gnd vdd FILL
XFILL_66_DFFSR_225 gnd vdd FILL
XFILL_9_BUFX4_105 gnd vdd FILL
XFILL_26_DFFSR_23 gnd vdd FILL
XFILL_66_DFFSR_236 gnd vdd FILL
XFILL_26_DFFSR_34 gnd vdd FILL
XFILL_66_DFFSR_247 gnd vdd FILL
XFILL_26_DFFSR_45 gnd vdd FILL
XFILL_26_DFFSR_56 gnd vdd FILL
XFILL_66_DFFSR_258 gnd vdd FILL
XFILL_66_DFFSR_269 gnd vdd FILL
XFILL_26_DFFSR_67 gnd vdd FILL
XFILL_26_DFFSR_78 gnd vdd FILL
XFILL_26_DFFSR_89 gnd vdd FILL
XFILL_66_DFFSR_11 gnd vdd FILL
XFILL_66_DFFSR_22 gnd vdd FILL
XFILL_66_DFFSR_33 gnd vdd FILL
XFILL_66_DFFSR_44 gnd vdd FILL
XFILL_1_MUX2X1_9 gnd vdd FILL
XFILL_66_DFFSR_55 gnd vdd FILL
XFILL_66_DFFSR_66 gnd vdd FILL
XFILL_66_DFFSR_77 gnd vdd FILL
XFILL_25_CLKBUF1_9 gnd vdd FILL
XFILL_7_4_0 gnd vdd FILL
XNAND3X1_10 AOI22X1_8/Y NAND3X1_10/B NOR3X1_42/Y gnd NOR3X1_43/A vdd NAND3X1
XNAND3X1_21 DFFSR_160/Q BUFX4_88/Y NOR2X1_36/Y gnd OAI21X1_29/C vdd NAND3X1
XFILL_66_DFFSR_88 gnd vdd FILL
XFILL_3_NOR2X1_19 gnd vdd FILL
XFILL_66_DFFSR_99 gnd vdd FILL
XNAND3X1_32 INVX1_137/A INVX1_134/Y INVX2_4/Y gnd OAI21X1_39/B vdd NAND3X1
XNAND3X1_43 NAND3X1_43/A NAND3X1_43/B OAI21X1_42/Y gnd NOR3X1_51/C vdd NAND3X1
XFILL_9_DFFSR_13 gnd vdd FILL
XFILL_4_BUFX4_1 gnd vdd FILL
XNAND3X1_54 NOR3X1_9/A DFFSR_199/D AND2X2_5/B gnd NOR3X1_4/B vdd NAND3X1
XFILL_29_DFFSR_9 gnd vdd FILL
XNAND3X1_65 NAND3X1_65/A NAND3X1_65/B NOR2X1_53/Y gnd NOR3X1_8/B vdd NAND3X1
XFILL_9_DFFSR_24 gnd vdd FILL
XFILL_7_NAND3X1_102 gnd vdd FILL
XFILL_9_DFFSR_35 gnd vdd FILL
XFILL_7_NAND3X1_113 gnd vdd FILL
XNAND3X1_76 DFFSR_103/Q BUFX4_2/Y NOR2X1_29/Y gnd OAI21X1_7/C vdd NAND3X1
XFILL_4_MUX2X1_180 gnd vdd FILL
XFILL_35_DFFSR_10 gnd vdd FILL
XFILL_35_DFFSR_21 gnd vdd FILL
XFILL_9_DFFSR_46 gnd vdd FILL
XNAND3X1_87 DFFSR_7/Q BUFX4_7/Y NOR3X1_9/Y gnd OAI21X1_10/C vdd NAND3X1
XFILL_7_NAND3X1_124 gnd vdd FILL
XFILL_4_MUX2X1_191 gnd vdd FILL
XFILL_9_DFFSR_57 gnd vdd FILL
XFILL_29_CLKBUF1_8 gnd vdd FILL
XFILL_35_DFFSR_32 gnd vdd FILL
XNOR2X1_10 NOR2X1_7/B NOR2X1_10/B gnd NOR2X1_12/B vdd NOR2X1
XNAND3X1_98 NOR2X1_28/A BUFX4_60/Y AND2X2_4/A gnd NAND3X1_98/Y vdd NAND3X1
XFILL_9_DFFSR_68 gnd vdd FILL
XNOR2X1_21 NOR2X1_21/A NOR2X1_21/B gnd INVX2_1/A vdd NOR2X1
XFILL_7_NOR2X1_18 gnd vdd FILL
XFILL_35_DFFSR_43 gnd vdd FILL
XNOR2X1_32 AND2X2_2/B AND2X2_2/A gnd BUFX4_8/A vdd NOR2X1
XFILL_9_DFFSR_79 gnd vdd FILL
XFILL_35_DFFSR_54 gnd vdd FILL
XNOR2X1_43 NOR3X1_49/B NOR2X1_52/B gnd NOR2X1_43/Y vdd NOR2X1
XFILL_7_NOR2X1_29 gnd vdd FILL
XFILL_35_DFFSR_65 gnd vdd FILL
XFILL_35_DFFSR_76 gnd vdd FILL
XNOR2X1_54 NOR3X1_51/Y AND2X2_5/Y gnd NOR2X1_54/Y vdd NOR2X1
XNOR2X1_65 INVX1_37/Y NOR2X1_80/B gnd NOR3X1_20/B vdd NOR2X1
XFILL_35_DFFSR_87 gnd vdd FILL
XNOR2X1_76 NOR2X1_76/A NOR2X1_76/B gnd NOR2X1_76/Y vdd NOR2X1
XFILL_35_DFFSR_98 gnd vdd FILL
XNOR2X1_87 INVX1_78/Y OAI22X1_1/D gnd NOR3X1_32/A vdd NOR2X1
XFILL_75_DFFSR_20 gnd vdd FILL
XNOR2X1_98 NOR2X1_98/A NOR2X1_98/B gnd NOR2X1_98/Y vdd NOR2X1
XFILL_75_DFFSR_31 gnd vdd FILL
XFILL_75_DFFSR_42 gnd vdd FILL
XFILL_15_3_0 gnd vdd FILL
XFILL_0_NOR2X1_109 gnd vdd FILL
XFILL_75_DFFSR_53 gnd vdd FILL
XFILL_75_DFFSR_64 gnd vdd FILL
XFILL_75_DFFSR_75 gnd vdd FILL
XFILL_75_DFFSR_86 gnd vdd FILL
XFILL_75_DFFSR_97 gnd vdd FILL
XFILL_3_INVX1_5 gnd vdd FILL
XFILL_10_NAND2X1_13 gnd vdd FILL
XFILL_10_NAND2X1_24 gnd vdd FILL
XFILL_10_NAND2X1_35 gnd vdd FILL
XFILL_10_NAND2X1_46 gnd vdd FILL
XFILL_10_NAND2X1_57 gnd vdd FILL
XFILL_44_DFFSR_30 gnd vdd FILL
XFILL_44_DFFSR_41 gnd vdd FILL
XFILL_15_NOR3X1_5 gnd vdd FILL
XFILL_8_OAI22X1_18 gnd vdd FILL
XFILL_44_DFFSR_52 gnd vdd FILL
XFILL_10_NAND2X1_68 gnd vdd FILL
XFILL_10_NAND2X1_79 gnd vdd FILL
XFILL_8_OAI22X1_29 gnd vdd FILL
XFILL_44_DFFSR_63 gnd vdd FILL
XFILL_44_DFFSR_74 gnd vdd FILL
XFILL_44_DFFSR_85 gnd vdd FILL
XFILL_82_DFFSR_190 gnd vdd FILL
XFILL_44_DFFSR_96 gnd vdd FILL
XFILL_33_DFFSR_203 gnd vdd FILL
XFILL_33_DFFSR_214 gnd vdd FILL
XFILL_33_DFFSR_225 gnd vdd FILL
XFILL_84_DFFSR_40 gnd vdd FILL
XFILL_84_DFFSR_51 gnd vdd FILL
XFILL_33_DFFSR_236 gnd vdd FILL
XFILL_7_NAND3X1_50 gnd vdd FILL
XFILL_33_DFFSR_247 gnd vdd FILL
XFILL_84_DFFSR_62 gnd vdd FILL
XFILL_2_DFFSR_260 gnd vdd FILL
XFILL_2_NAND3X1_120 gnd vdd FILL
XFILL_2_DFFSR_271 gnd vdd FILL
XFILL_7_NAND3X1_61 gnd vdd FILL
XFILL_33_DFFSR_258 gnd vdd FILL
XFILL_4_INVX4_1 gnd vdd FILL
XFILL_2_NAND3X1_131 gnd vdd FILL
XFILL_33_DFFSR_269 gnd vdd FILL
XFILL_84_DFFSR_73 gnd vdd FILL
XFILL_84_DFFSR_84 gnd vdd FILL
XFILL_13_DFFSR_40 gnd vdd FILL
XFILL_7_NAND3X1_72 gnd vdd FILL
XFILL_84_DFFSR_95 gnd vdd FILL
XFILL_13_DFFSR_51 gnd vdd FILL
XFILL_60_DFFSR_103 gnd vdd FILL
XFILL_7_NAND3X1_83 gnd vdd FILL
XFILL_37_DFFSR_202 gnd vdd FILL
XFILL_7_NAND3X1_94 gnd vdd FILL
XFILL_13_DFFSR_62 gnd vdd FILL
XFILL_37_DFFSR_213 gnd vdd FILL
XFILL_60_DFFSR_114 gnd vdd FILL
XFILL_13_DFFSR_73 gnd vdd FILL
XFILL_37_DFFSR_224 gnd vdd FILL
XFILL_60_DFFSR_125 gnd vdd FILL
XFILL_60_DFFSR_136 gnd vdd FILL
XFILL_13_DFFSR_84 gnd vdd FILL
XFILL_37_DFFSR_235 gnd vdd FILL
XFILL_13_DFFSR_95 gnd vdd FILL
XFILL_60_DFFSR_147 gnd vdd FILL
XFILL_60_DFFSR_158 gnd vdd FILL
XFILL_37_DFFSR_246 gnd vdd FILL
XFILL_6_DFFSR_270 gnd vdd FILL
XFILL_37_DFFSR_257 gnd vdd FILL
XFILL_37_DFFSR_268 gnd vdd FILL
XFILL_60_DFFSR_169 gnd vdd FILL
XFILL_3_MUX2X1_15 gnd vdd FILL
XNAND2X1_9 INVX2_1/A NOR2X1_24/Y gnd NAND2X1_9/Y vdd NAND2X1
XFILL_24_NOR3X1_3 gnd vdd FILL
XFILL_64_DFFSR_102 gnd vdd FILL
XFILL_10_AOI22X1_11 gnd vdd FILL
XFILL_3_MUX2X1_26 gnd vdd FILL
XFILL_53_DFFSR_50 gnd vdd FILL
XFILL_19_CLKBUF1_16 gnd vdd FILL
XFILL_3_MUX2X1_37 gnd vdd FILL
XFILL_64_DFFSR_113 gnd vdd FILL
XFILL_53_DFFSR_61 gnd vdd FILL
XFILL_66_7_1 gnd vdd FILL
XFILL_3_MUX2X1_48 gnd vdd FILL
XFILL_53_DFFSR_72 gnd vdd FILL
XFILL_64_DFFSR_124 gnd vdd FILL
XFILL_3_MUX2X1_59 gnd vdd FILL
XFILL_19_CLKBUF1_27 gnd vdd FILL
XFILL_53_DFFSR_83 gnd vdd FILL
XFILL_19_CLKBUF1_38 gnd vdd FILL
XFILL_64_DFFSR_135 gnd vdd FILL
XFILL_65_2_0 gnd vdd FILL
XFILL_64_DFFSR_146 gnd vdd FILL
XFILL_14_AOI21X1_13 gnd vdd FILL
XFILL_53_DFFSR_94 gnd vdd FILL
XFILL_64_DFFSR_157 gnd vdd FILL
XFILL_14_AOI21X1_24 gnd vdd FILL
XFILL_64_DFFSR_168 gnd vdd FILL
XFILL_7_MUX2X1_14 gnd vdd FILL
XFILL_14_AOI21X1_35 gnd vdd FILL
XFILL_0_NAND2X1_30 gnd vdd FILL
XFILL_14_AOI21X1_46 gnd vdd FILL
XFILL_64_DFFSR_179 gnd vdd FILL
XNOR2X1_100 OAI22X1_39/Y OAI22X1_40/Y gnd NOR2X1_100/Y vdd NOR2X1
XFILL_7_MUX2X1_25 gnd vdd FILL
XFILL_68_DFFSR_101 gnd vdd FILL
XFILL_0_NAND2X1_41 gnd vdd FILL
XNOR2X1_111 INVX1_133/A INVX1_131/Y gnd OAI21X1_1/A vdd NOR2X1
XFILL_14_AOI21X1_57 gnd vdd FILL
XFILL_0_NAND2X1_52 gnd vdd FILL
XFILL_7_MUX2X1_36 gnd vdd FILL
XFILL_68_DFFSR_112 gnd vdd FILL
XMUX2X1_50 INVX1_63/Y BUFX4_85/Y NAND2X1_8/Y gnd MUX2X1_50/Y vdd MUX2X1
XFILL_14_AOI21X1_68 gnd vdd FILL
XFILL_0_NAND2X1_63 gnd vdd FILL
XFILL_7_MUX2X1_47 gnd vdd FILL
XMUX2X1_61 MUX2X1_6/B INVX1_74/Y NOR2X1_22/Y gnd MUX2X1_61/Y vdd MUX2X1
XNOR2X1_122 BUFX2_7/A INVX2_3/Y gnd NOR2X1_122/Y vdd NOR2X1
XFILL_68_DFFSR_123 gnd vdd FILL
XFILL_0_NAND2X1_74 gnd vdd FILL
XNOR2X1_133 DFFSR_141/Q AOI21X1_7/B gnd AOI21X1_6/C vdd NOR2X1
XFILL_7_MUX2X1_58 gnd vdd FILL
XFILL_14_AOI21X1_79 gnd vdd FILL
XMUX2X1_72 INVX1_85/Y BUFX4_86/Y OR2X2_1/Y gnd MUX2X1_72/Y vdd MUX2X1
XFILL_68_DFFSR_134 gnd vdd FILL
XFILL_7_MUX2X1_69 gnd vdd FILL
XMUX2X1_83 INVX1_96/Y MUX2X1_8/A MUX2X1_86/S gnd MUX2X1_83/Y vdd MUX2X1
XNOR2X1_144 DFFSR_103/Q AOI21X1_9/B gnd AOI21X1_8/C vdd NOR2X1
XFILL_0_NAND2X1_85 gnd vdd FILL
XFILL_11_OAI21X1_2 gnd vdd FILL
XFILL_68_DFFSR_145 gnd vdd FILL
XNOR2X1_155 NOR2X1_57/A NAND2X1_3/Y gnd NOR2X1_155/Y vdd NOR2X1
XFILL_68_DFFSR_156 gnd vdd FILL
XMUX2X1_94 MUX2X1_94/A BUFX4_75/Y MUX2X1_95/S gnd MUX2X1_94/Y vdd MUX2X1
XFILL_22_DFFSR_60 gnd vdd FILL
XFILL_0_NAND2X1_96 gnd vdd FILL
XNOR2X1_166 NOR2X1_7/A NAND2X1_3/Y gnd NOR2X1_166/Y vdd NOR2X1
XFILL_68_DFFSR_167 gnd vdd FILL
XFILL_22_DFFSR_71 gnd vdd FILL
XFILL_22_DFFSR_82 gnd vdd FILL
XNOR2X1_177 NOR2X1_7/B INVX1_68/Y gnd NOR2X1_181/B vdd NOR2X1
XFILL_68_DFFSR_178 gnd vdd FILL
XNOR2X1_188 DFFSR_20/Q NOR2X1_190/B gnd NOR2X1_188/Y vdd NOR2X1
XFILL_22_DFFSR_93 gnd vdd FILL
XNOR2X1_199 DFFSR_6/Q NOR2X1_202/B gnd NOR2X1_199/Y vdd NOR2X1
XFILL_68_DFFSR_189 gnd vdd FILL
XFILL_7_NOR3X1_4 gnd vdd FILL
XFILL_15_OAI21X1_1 gnd vdd FILL
XFILL_62_DFFSR_70 gnd vdd FILL
XFILL_62_DFFSR_81 gnd vdd FILL
XFILL_62_DFFSR_92 gnd vdd FILL
XFILL_26_CLKBUF1_40 gnd vdd FILL
XFILL_46_DFFSR_3 gnd vdd FILL
XFILL_5_DFFSR_50 gnd vdd FILL
XMUX2X1_106 BUFX4_81/Y OAI22X1_4/A MUX2X1_1/S gnd DFFSR_183/D vdd MUX2X1
XFILL_5_DFFSR_61 gnd vdd FILL
XMUX2X1_117 INVX1_159/Y BUFX4_81/Y NAND2X1_78/Y gnd DFFSR_134/D vdd MUX2X1
XFILL_9_CLKBUF1_11 gnd vdd FILL
XFILL_5_DFFSR_72 gnd vdd FILL
XFILL_5_DFFSR_83 gnd vdd FILL
XFILL_9_CLKBUF1_22 gnd vdd FILL
XFILL_23_MUX2X1_12 gnd vdd FILL
XFILL_9_CLKBUF1_33 gnd vdd FILL
XMUX2X1_128 INVX1_172/Y BUFX4_77/Y NAND2X1_89/Y gnd DFFSR_128/D vdd MUX2X1
XFILL_23_MUX2X1_23 gnd vdd FILL
XMUX2X1_139 INVX1_183/Y MUX2X1_4/B NAND3X1_1/Y gnd DFFSR_111/D vdd MUX2X1
XFILL_5_DFFSR_94 gnd vdd FILL
XFILL_31_DFFSR_80 gnd vdd FILL
XFILL_23_MUX2X1_34 gnd vdd FILL
XFILL_17_MUX2X1_107 gnd vdd FILL
XFILL_31_DFFSR_91 gnd vdd FILL
XFILL_23_MUX2X1_45 gnd vdd FILL
XFILL_4_AOI21X1_30 gnd vdd FILL
XFILL_17_MUX2X1_118 gnd vdd FILL
XFILL_23_MUX2X1_56 gnd vdd FILL
XFILL_17_MUX2X1_129 gnd vdd FILL
XFILL_23_MUX2X1_67 gnd vdd FILL
XFILL_4_AOI21X1_41 gnd vdd FILL
XFILL_23_MUX2X1_78 gnd vdd FILL
XFILL_4_AOI21X1_52 gnd vdd FILL
XFILL_14_OAI22X1_10 gnd vdd FILL
XFILL_23_MUX2X1_89 gnd vdd FILL
XFILL_4_AOI21X1_63 gnd vdd FILL
XFILL_9_BUFX2_8 gnd vdd FILL
XFILL_4_AOI21X1_74 gnd vdd FILL
XFILL_14_OAI22X1_21 gnd vdd FILL
XFILL_14_OAI22X1_32 gnd vdd FILL
XFILL_14_OAI22X1_43 gnd vdd FILL
XINVX1_13 INVX1_13/A gnd INVX1_13/Y vdd INVX1
XINVX1_24 INVX1_24/A gnd INVX1_24/Y vdd INVX1
XFILL_71_DFFSR_90 gnd vdd FILL
XINVX1_35 INVX1_35/A gnd MUX2X1_2/B vdd INVX1
XINVX1_46 INVX1_46/A gnd INVX1_46/Y vdd INVX1
XFILL_30_DFFSR_9 gnd vdd FILL
XFILL_7_NOR2X1_140 gnd vdd FILL
XINVX1_57 INVX1_57/A gnd INVX1_57/Y vdd INVX1
XFILL_7_NOR2X1_151 gnd vdd FILL
XINVX1_68 INVX1_68/A gnd INVX1_68/Y vdd INVX1
XFILL_57_7_1 gnd vdd FILL
XFILL_7_NOR2X1_162 gnd vdd FILL
XINVX1_79 INVX1_79/A gnd INVX1_79/Y vdd INVX1
XFILL_7_NOR2X1_173 gnd vdd FILL
XFILL_31_DFFSR_102 gnd vdd FILL
XFILL_56_2_0 gnd vdd FILL
XFILL_7_NOR2X1_184 gnd vdd FILL
XFILL_7_NOR2X1_195 gnd vdd FILL
XFILL_31_DFFSR_113 gnd vdd FILL
XFILL_68_DFFSR_7 gnd vdd FILL
XFILL_31_DFFSR_124 gnd vdd FILL
XFILL_31_DFFSR_135 gnd vdd FILL
XFILL_31_DFFSR_146 gnd vdd FILL
XFILL_11_NOR2X1_201 gnd vdd FILL
XFILL_31_DFFSR_157 gnd vdd FILL
XFILL_0_DFFSR_170 gnd vdd FILL
XFILL_31_DFFSR_168 gnd vdd FILL
XFILL_0_DFFSR_181 gnd vdd FILL
XFILL_31_DFFSR_179 gnd vdd FILL
XFILL_0_DFFSR_192 gnd vdd FILL
XFILL_35_DFFSR_101 gnd vdd FILL
XFILL_35_DFFSR_112 gnd vdd FILL
XFILL_35_DFFSR_123 gnd vdd FILL
XFILL_35_DFFSR_134 gnd vdd FILL
XFILL_35_DFFSR_145 gnd vdd FILL
XFILL_35_DFFSR_156 gnd vdd FILL
XFILL_35_DFFSR_167 gnd vdd FILL
XFILL_4_DFFSR_180 gnd vdd FILL
XFILL_40_6_1 gnd vdd FILL
XFILL_35_DFFSR_178 gnd vdd FILL
XFILL_4_DFFSR_191 gnd vdd FILL
XFILL_7_MUX2X1_102 gnd vdd FILL
XFILL_39_DFFSR_100 gnd vdd FILL
XFILL_35_DFFSR_189 gnd vdd FILL
XFILL_7_MUX2X1_113 gnd vdd FILL
XFILL_39_DFFSR_111 gnd vdd FILL
XFILL_7_MUX2X1_124 gnd vdd FILL
XFILL_39_DFFSR_122 gnd vdd FILL
XFILL_7_MUX2X1_135 gnd vdd FILL
XFILL_39_DFFSR_133 gnd vdd FILL
XFILL_7_MUX2X1_146 gnd vdd FILL
XFILL_39_DFFSR_144 gnd vdd FILL
XFILL_8_BUFX4_2 gnd vdd FILL
XFILL_39_DFFSR_155 gnd vdd FILL
XFILL_7_MUX2X1_157 gnd vdd FILL
XFILL_7_MUX2X1_168 gnd vdd FILL
XFILL_39_DFFSR_166 gnd vdd FILL
XFILL_39_DFFSR_177 gnd vdd FILL
XFILL_7_MUX2X1_179 gnd vdd FILL
XFILL_31_NOR3X1_13 gnd vdd FILL
XFILL_8_DFFSR_190 gnd vdd FILL
XFILL_31_NOR3X1_24 gnd vdd FILL
XFILL_39_DFFSR_188 gnd vdd FILL
XFILL_31_NOR3X1_35 gnd vdd FILL
XFILL_39_DFFSR_199 gnd vdd FILL
XFILL_81_DFFSR_202 gnd vdd FILL
XFILL_31_NOR3X1_46 gnd vdd FILL
XFILL_81_DFFSR_213 gnd vdd FILL
XFILL_8_OAI21X1_40 gnd vdd FILL
XFILL_81_DFFSR_224 gnd vdd FILL
XFILL_81_DFFSR_235 gnd vdd FILL
XFILL_81_DFFSR_246 gnd vdd FILL
XFILL_81_DFFSR_257 gnd vdd FILL
XFILL_81_DFFSR_268 gnd vdd FILL
XFILL_85_DFFSR_201 gnd vdd FILL
XFILL_85_DFFSR_212 gnd vdd FILL
XFILL_85_DFFSR_223 gnd vdd FILL
XFILL_85_DFFSR_234 gnd vdd FILL
XFILL_12_AOI21X1_8 gnd vdd FILL
XFILL_7_INVX1_6 gnd vdd FILL
XFILL_85_DFFSR_245 gnd vdd FILL
XFILL_85_DFFSR_256 gnd vdd FILL
XFILL_85_DFFSR_267 gnd vdd FILL
XFILL_66_9 gnd vdd FILL
XFILL_48_7_1 gnd vdd FILL
XFILL_1_INVX1_140 gnd vdd FILL
XFILL_1_INVX1_151 gnd vdd FILL
XFILL_1_INVX1_162 gnd vdd FILL
XFILL_47_2_0 gnd vdd FILL
XFILL_8_NAND3X1_103 gnd vdd FILL
XFILL_1_INVX1_173 gnd vdd FILL
XFILL_8_NAND3X1_114 gnd vdd FILL
XFILL_1_INVX1_184 gnd vdd FILL
XFILL_8_NAND3X1_125 gnd vdd FILL
XFILL_1_INVX1_195 gnd vdd FILL
XFILL_5_INVX1_150 gnd vdd FILL
XFILL_5_INVX1_161 gnd vdd FILL
XFILL_5_INVX1_172 gnd vdd FILL
XFILL_5_INVX1_183 gnd vdd FILL
XFILL_5_INVX1_194 gnd vdd FILL
XFILL_31_6_1 gnd vdd FILL
XFILL_30_1_0 gnd vdd FILL
XFILL_3_OAI22X1_1 gnd vdd FILL
XFILL_3_NAND2X1_18 gnd vdd FILL
XFILL_3_NAND2X1_29 gnd vdd FILL
XFILL_85_DFFSR_1 gnd vdd FILL
XFILL_0_AND2X2_8 gnd vdd FILL
XFILL_3_NAND3X1_110 gnd vdd FILL
XFILL_3_NAND3X1_121 gnd vdd FILL
XFILL_45_DFFSR_19 gnd vdd FILL
XFILL_13_MUX2X1_160 gnd vdd FILL
XFILL_3_NAND3X1_132 gnd vdd FILL
XFILL_13_MUX2X1_171 gnd vdd FILL
XFILL_13_MUX2X1_182 gnd vdd FILL
XFILL_52_DFFSR_201 gnd vdd FILL
XFILL_13_MUX2X1_193 gnd vdd FILL
XFILL_52_DFFSR_212 gnd vdd FILL
XFILL_52_DFFSR_223 gnd vdd FILL
XFILL_52_DFFSR_234 gnd vdd FILL
XFILL_52_DFFSR_245 gnd vdd FILL
XFILL_39_7_1 gnd vdd FILL
XFILL_85_DFFSR_18 gnd vdd FILL
XFILL_52_DFFSR_256 gnd vdd FILL
XFILL_52_DFFSR_267 gnd vdd FILL
XFILL_85_DFFSR_29 gnd vdd FILL
XFILL_12_DFFSR_6 gnd vdd FILL
XFILL_38_2_0 gnd vdd FILL
XFILL_56_DFFSR_200 gnd vdd FILL
XFILL_29_CLKBUF1_17 gnd vdd FILL
XFILL_56_DFFSR_211 gnd vdd FILL
XFILL_14_DFFSR_18 gnd vdd FILL
XFILL_29_CLKBUF1_28 gnd vdd FILL
XFILL_56_DFFSR_222 gnd vdd FILL
XFILL_14_DFFSR_29 gnd vdd FILL
XFILL_56_DFFSR_233 gnd vdd FILL
XFILL_29_CLKBUF1_39 gnd vdd FILL
XFILL_56_DFFSR_244 gnd vdd FILL
XFILL_56_DFFSR_255 gnd vdd FILL
XFILL_56_DFFSR_266 gnd vdd FILL
XFILL_11_CLKBUF1_7 gnd vdd FILL
XFILL_83_DFFSR_100 gnd vdd FILL
XFILL_83_DFFSR_111 gnd vdd FILL
XFILL_54_DFFSR_17 gnd vdd FILL
XFILL_7_AOI21X1_18 gnd vdd FILL
XOAI22X1_19 INVX1_87/Y OAI22X1_8/B INVX1_98/Y OAI22X1_8/D gnd NOR3X1_28/A vdd OAI22X1
XFILL_54_DFFSR_28 gnd vdd FILL
XFILL_83_DFFSR_122 gnd vdd FILL
XFILL_83_DFFSR_133 gnd vdd FILL
XFILL_7_AOI21X1_29 gnd vdd FILL
XFILL_54_DFFSR_39 gnd vdd FILL
XFILL_83_DFFSR_144 gnd vdd FILL
XFILL_83_DFFSR_155 gnd vdd FILL
XFILL_83_DFFSR_166 gnd vdd FILL
XFILL_22_6_1 gnd vdd FILL
XFILL_83_DFFSR_177 gnd vdd FILL
XFILL_15_CLKBUF1_6 gnd vdd FILL
XFILL_83_DFFSR_188 gnd vdd FILL
XFILL_3_DFFSR_203 gnd vdd FILL
XFILL_0_NAND3X1_3 gnd vdd FILL
XFILL_87_DFFSR_110 gnd vdd FILL
XFILL_83_DFFSR_199 gnd vdd FILL
XFILL_21_1_0 gnd vdd FILL
XFILL_3_DFFSR_214 gnd vdd FILL
XFILL_87_DFFSR_121 gnd vdd FILL
XFILL_3_DFFSR_225 gnd vdd FILL
XFILL_87_DFFSR_132 gnd vdd FILL
XFILL_3_DFFSR_236 gnd vdd FILL
XFILL_87_DFFSR_143 gnd vdd FILL
XFILL_3_DFFSR_247 gnd vdd FILL
XFILL_87_DFFSR_154 gnd vdd FILL
XFILL_11_BUFX4_101 gnd vdd FILL
XFILL_23_DFFSR_16 gnd vdd FILL
XFILL_3_DFFSR_258 gnd vdd FILL
XFILL_3_DFFSR_269 gnd vdd FILL
XFILL_87_DFFSR_165 gnd vdd FILL
XFILL_23_DFFSR_27 gnd vdd FILL
XFILL_87_DFFSR_176 gnd vdd FILL
XFILL_23_DFFSR_38 gnd vdd FILL
XFILL_19_CLKBUF1_5 gnd vdd FILL
XFILL_7_DFFSR_202 gnd vdd FILL
XFILL_14_BUFX4_70 gnd vdd FILL
XFILL_87_DFFSR_187 gnd vdd FILL
XFILL_23_DFFSR_49 gnd vdd FILL
XFILL_4_NAND3X1_2 gnd vdd FILL
XFILL_14_BUFX4_81 gnd vdd FILL
XFILL_7_DFFSR_213 gnd vdd FILL
XFILL_87_DFFSR_198 gnd vdd FILL
XFILL_14_BUFX4_92 gnd vdd FILL
XFILL_7_DFFSR_224 gnd vdd FILL
XFILL_7_DFFSR_235 gnd vdd FILL
XDFFSR_260 INVX1_42/A DFFSR_9/CLK DFFSR_9/R vdd MUX2X1_29/Y gnd vdd DFFSR
XFILL_7_DFFSR_246 gnd vdd FILL
XDFFSR_271 NOR2X1_3/A DFFSR_6/CLK DFFSR_6/R vdd DFFSR_271/D gnd vdd DFFSR
XFILL_63_DFFSR_15 gnd vdd FILL
XFILL_7_DFFSR_257 gnd vdd FILL
XFILL_15_BUFX4_100 gnd vdd FILL
XFILL_7_DFFSR_268 gnd vdd FILL
XFILL_63_DFFSR_26 gnd vdd FILL
XFILL_63_DFFSR_37 gnd vdd FILL
XFILL_63_DFFSR_48 gnd vdd FILL
XFILL_8_NAND3X1_1 gnd vdd FILL
XFILL_63_DFFSR_59 gnd vdd FILL
XFILL_6_DFFSR_17 gnd vdd FILL
XFILL_6_DFFSR_28 gnd vdd FILL
XFILL_32_DFFSR_14 gnd vdd FILL
XFILL_6_DFFSR_39 gnd vdd FILL
XFILL_32_DFFSR_25 gnd vdd FILL
XFILL_32_DFFSR_36 gnd vdd FILL
XFILL_5_7_1 gnd vdd FILL
XFILL_0_AOI22X1_8 gnd vdd FILL
XFILL_32_DFFSR_47 gnd vdd FILL
XFILL_32_DFFSR_58 gnd vdd FILL
XFILL_7_OAI22X1_15 gnd vdd FILL
XFILL_4_2_0 gnd vdd FILL
XFILL_32_DFFSR_69 gnd vdd FILL
XFILL_7_OAI22X1_26 gnd vdd FILL
XFILL_29_2_0 gnd vdd FILL
XFILL_7_OAI22X1_37 gnd vdd FILL
XFILL_7_OAI22X1_48 gnd vdd FILL
XFILL_72_DFFSR_13 gnd vdd FILL
XFILL_0_INVX1_207 gnd vdd FILL
XFILL_23_DFFSR_200 gnd vdd FILL
XFILL_72_DFFSR_24 gnd vdd FILL
XFILL_0_INVX1_218 gnd vdd FILL
XFILL_23_DFFSR_211 gnd vdd FILL
XFILL_72_DFFSR_35 gnd vdd FILL
XFILL_23_DFFSR_222 gnd vdd FILL
XFILL_72_DFFSR_46 gnd vdd FILL
XFILL_23_DFFSR_233 gnd vdd FILL
XFILL_15_MUX2X1_3 gnd vdd FILL
XFILL_4_AOI22X1_7 gnd vdd FILL
XFILL_72_DFFSR_57 gnd vdd FILL
XFILL_72_DFFSR_68 gnd vdd FILL
XFILL_23_DFFSR_244 gnd vdd FILL
XFILL_23_DFFSR_255 gnd vdd FILL
XFILL_72_DFFSR_79 gnd vdd FILL
XFILL_23_DFFSR_266 gnd vdd FILL
XFILL_4_INVX1_206 gnd vdd FILL
XFILL_50_DFFSR_100 gnd vdd FILL
XFILL_6_NAND3X1_80 gnd vdd FILL
XFILL_6_NAND3X1_91 gnd vdd FILL
XFILL_50_DFFSR_111 gnd vdd FILL
XFILL_4_INVX1_217 gnd vdd FILL
XFILL_27_DFFSR_210 gnd vdd FILL
XFILL_4_INVX1_228 gnd vdd FILL
XFILL_4_NOR2X1_206 gnd vdd FILL
XFILL_13_6_1 gnd vdd FILL
XFILL_27_DFFSR_221 gnd vdd FILL
XFILL_50_DFFSR_122 gnd vdd FILL
XFILL_8_AOI22X1_6 gnd vdd FILL
XFILL_50_DFFSR_133 gnd vdd FILL
XFILL_27_DFFSR_232 gnd vdd FILL
XFILL_27_DFFSR_243 gnd vdd FILL
XFILL_50_DFFSR_144 gnd vdd FILL
XFILL_41_DFFSR_12 gnd vdd FILL
XFILL_50_DFFSR_155 gnd vdd FILL
XFILL_12_1_0 gnd vdd FILL
XFILL_41_DFFSR_23 gnd vdd FILL
XFILL_6_BUFX4_80 gnd vdd FILL
XFILL_27_DFFSR_254 gnd vdd FILL
XFILL_41_DFFSR_34 gnd vdd FILL
XFILL_6_BUFX4_91 gnd vdd FILL
XFILL_12_NOR3X1_9 gnd vdd FILL
XFILL_41_DFFSR_45 gnd vdd FILL
XFILL_50_DFFSR_166 gnd vdd FILL
XFILL_27_DFFSR_265 gnd vdd FILL
XFILL_41_DFFSR_56 gnd vdd FILL
XFILL_50_DFFSR_177 gnd vdd FILL
XFILL_0_OAI21X1_17 gnd vdd FILL
XFILL_50_DFFSR_188 gnd vdd FILL
XFILL_0_OAI21X1_28 gnd vdd FILL
XFILL_41_DFFSR_67 gnd vdd FILL
XFILL_54_DFFSR_110 gnd vdd FILL
XFILL_50_DFFSR_199 gnd vdd FILL
XFILL_18_CLKBUF1_13 gnd vdd FILL
XFILL_41_DFFSR_78 gnd vdd FILL
XFILL_18_CLKBUF1_24 gnd vdd FILL
XFILL_54_DFFSR_121 gnd vdd FILL
XFILL_0_OAI21X1_39 gnd vdd FILL
XFILL_41_DFFSR_89 gnd vdd FILL
XFILL_54_DFFSR_132 gnd vdd FILL
XFILL_81_DFFSR_11 gnd vdd FILL
XFILL_18_CLKBUF1_35 gnd vdd FILL
XFILL_54_DFFSR_143 gnd vdd FILL
XFILL_13_AOI21X1_10 gnd vdd FILL
XFILL_54_DFFSR_154 gnd vdd FILL
XFILL_13_AOI21X1_21 gnd vdd FILL
XFILL_81_DFFSR_22 gnd vdd FILL
XFILL_54_DFFSR_165 gnd vdd FILL
XFILL_81_DFFSR_33 gnd vdd FILL
XFILL_13_AOI21X1_32 gnd vdd FILL
XFILL_81_DFFSR_44 gnd vdd FILL
XFILL_13_AOI21X1_43 gnd vdd FILL
XFILL_81_DFFSR_55 gnd vdd FILL
XFILL_10_DFFSR_11 gnd vdd FILL
XFILL_54_DFFSR_176 gnd vdd FILL
XFILL_54_DFFSR_187 gnd vdd FILL
XFILL_13_AOI21X1_54 gnd vdd FILL
XFILL_81_DFFSR_66 gnd vdd FILL
XFILL_54_DFFSR_198 gnd vdd FILL
XFILL_10_DFFSR_22 gnd vdd FILL
XFILL_13_AOI21X1_65 gnd vdd FILL
XFILL_81_DFFSR_77 gnd vdd FILL
XFILL_58_DFFSR_120 gnd vdd FILL
XFILL_10_DFFSR_33 gnd vdd FILL
XFILL_81_DFFSR_88 gnd vdd FILL
XFILL_13_AOI21X1_76 gnd vdd FILL
XFILL_10_DFFSR_44 gnd vdd FILL
XFILL_58_DFFSR_131 gnd vdd FILL
XFILL_10_DFFSR_55 gnd vdd FILL
XFILL_81_DFFSR_99 gnd vdd FILL
XFILL_58_DFFSR_142 gnd vdd FILL
XFILL_10_DFFSR_66 gnd vdd FILL
XFILL_58_DFFSR_153 gnd vdd FILL
XFILL_8_NOR2X1_4 gnd vdd FILL
XFILL_10_DFFSR_77 gnd vdd FILL
XFILL_58_DFFSR_164 gnd vdd FILL
XFILL_58_DFFSR_175 gnd vdd FILL
XFILL_10_DFFSR_88 gnd vdd FILL
XFILL_1_DFFSR_102 gnd vdd FILL
XFILL_10_DFFSR_99 gnd vdd FILL
XFILL_50_DFFSR_10 gnd vdd FILL
XFILL_50_DFFSR_21 gnd vdd FILL
XFILL_58_DFFSR_186 gnd vdd FILL
XFILL_1_DFFSR_113 gnd vdd FILL
XFILL_58_DFFSR_197 gnd vdd FILL
XFILL_1_DFFSR_124 gnd vdd FILL
XFILL_50_DFFSR_32 gnd vdd FILL
XFILL_50_DFFSR_43 gnd vdd FILL
XFILL_1_DFFSR_135 gnd vdd FILL
XFILL_8_4 gnd vdd FILL
XFILL_21_NOR3X1_7 gnd vdd FILL
XFILL_1_DFFSR_146 gnd vdd FILL
XFILL_50_DFFSR_54 gnd vdd FILL
XFILL_1_DFFSR_157 gnd vdd FILL
XFILL_50_DFFSR_65 gnd vdd FILL
XFILL_50_DFFSR_76 gnd vdd FILL
XFILL_1_DFFSR_168 gnd vdd FILL
XFILL_1_DFFSR_179 gnd vdd FILL
XFILL_50_DFFSR_87 gnd vdd FILL
XFILL_50_DFFSR_98 gnd vdd FILL
XFILL_5_DFFSR_101 gnd vdd FILL
XFILL_5_DFFSR_112 gnd vdd FILL
XFILL_7_MUX2X1_2 gnd vdd FILL
XFILL_5_DFFSR_123 gnd vdd FILL
XFILL_5_DFFSR_134 gnd vdd FILL
XFILL_57_5 gnd vdd FILL
XFILL_5_DFFSR_145 gnd vdd FILL
XFILL_5_DFFSR_156 gnd vdd FILL
XFILL_51_DFFSR_4 gnd vdd FILL
XFILL_5_DFFSR_167 gnd vdd FILL
XFILL_5_DFFSR_178 gnd vdd FILL
XFILL_9_NAND3X1_104 gnd vdd FILL
XFILL_63_5_1 gnd vdd FILL
XFILL_9_DFFSR_100 gnd vdd FILL
XFILL_9_NAND3X1_115 gnd vdd FILL
XFILL_5_DFFSR_189 gnd vdd FILL
XFILL_9_DFFSR_111 gnd vdd FILL
XFILL_9_NAND3X1_126 gnd vdd FILL
XFILL_8_CLKBUF1_30 gnd vdd FILL
XFILL_9_DFFSR_122 gnd vdd FILL
XFILL_13_MUX2X1_20 gnd vdd FILL
XFILL_8_CLKBUF1_41 gnd vdd FILL
XFILL_62_0_0 gnd vdd FILL
XFILL_9_DFFSR_133 gnd vdd FILL
XFILL_16_MUX2X1_104 gnd vdd FILL
XFILL_13_MUX2X1_31 gnd vdd FILL
XFILL_9_DFFSR_144 gnd vdd FILL
XFILL_16_MUX2X1_115 gnd vdd FILL
XFILL_13_MUX2X1_42 gnd vdd FILL
XFILL_4_NOR3X1_8 gnd vdd FILL
XFILL_13_MUX2X1_53 gnd vdd FILL
XFILL_9_DFFSR_155 gnd vdd FILL
XFILL_13_MUX2X1_64 gnd vdd FILL
XFILL_16_MUX2X1_126 gnd vdd FILL
XFILL_9_DFFSR_166 gnd vdd FILL
XFILL_9_DFFSR_177 gnd vdd FILL
XFILL_13_MUX2X1_75 gnd vdd FILL
XFILL_16_MUX2X1_137 gnd vdd FILL
XFILL_30_NOR3X1_5 gnd vdd FILL
XFILL_1_NOR3X1_13 gnd vdd FILL
XFILL_16_MUX2X1_148 gnd vdd FILL
XFILL_13_MUX2X1_86 gnd vdd FILL
XFILL_1_NOR3X1_24 gnd vdd FILL
XFILL_16_MUX2X1_159 gnd vdd FILL
XFILL_9_DFFSR_188 gnd vdd FILL
XFILL_3_AOI21X1_60 gnd vdd FILL
XFILL_13_MUX2X1_97 gnd vdd FILL
XFILL_3_AOI21X1_71 gnd vdd FILL
XFILL_1_NOR3X1_35 gnd vdd FILL
XFILL_9_DFFSR_199 gnd vdd FILL
XOAI21X1_30 INVX1_210/Y OAI21X1_5/B OAI21X1_30/C gnd OAI21X1_30/Y vdd OAI21X1
XFILL_1_NOR3X1_46 gnd vdd FILL
XFILL_17_MUX2X1_30 gnd vdd FILL
XOAI21X1_41 OAI21X1_41/A AOI22X1_3/A INVX2_4/Y gnd OAI21X1_41/Y vdd OAI21X1
XFILL_13_OAI22X1_40 gnd vdd FILL
XFILL_13_OAI22X1_51 gnd vdd FILL
XFILL_17_MUX2X1_41 gnd vdd FILL
XFILL_17_MUX2X1_52 gnd vdd FILL
XFILL_17_MUX2X1_63 gnd vdd FILL
XFILL_2_DFFSR_10 gnd vdd FILL
XFILL_2_DFFSR_21 gnd vdd FILL
XFILL_17_MUX2X1_74 gnd vdd FILL
XFILL_3_DFFSR_9 gnd vdd FILL
XFILL_5_NOR3X1_12 gnd vdd FILL
XFILL_2_DFFSR_32 gnd vdd FILL
XFILL_17_MUX2X1_85 gnd vdd FILL
XFILL_5_NOR3X1_23 gnd vdd FILL
XFILL_5_NOR3X1_34 gnd vdd FILL
XFILL_2_DFFSR_43 gnd vdd FILL
XFILL_17_MUX2X1_96 gnd vdd FILL
XFILL_6_NOR2X1_170 gnd vdd FILL
XFILL_16_DFFSR_7 gnd vdd FILL
XFILL_6_NOR2X1_181 gnd vdd FILL
XFILL_2_DFFSR_54 gnd vdd FILL
XFILL_5_NOR3X1_45 gnd vdd FILL
XFILL_73_DFFSR_8 gnd vdd FILL
XFILL_2_DFFSR_65 gnd vdd FILL
XFILL_21_DFFSR_110 gnd vdd FILL
XFILL_2_DFFSR_76 gnd vdd FILL
XFILL_6_NOR2X1_192 gnd vdd FILL
XFILL_2_DFFSR_87 gnd vdd FILL
XFILL_21_DFFSR_121 gnd vdd FILL
XFILL_21_DFFSR_132 gnd vdd FILL
XFILL_21_DFFSR_143 gnd vdd FILL
XFILL_2_DFFSR_98 gnd vdd FILL
XFILL_21_DFFSR_154 gnd vdd FILL
XFILL_9_NOR3X1_11 gnd vdd FILL
XFILL_21_DFFSR_165 gnd vdd FILL
XFILL_9_NOR3X1_22 gnd vdd FILL
XFILL_2_INVX1_105 gnd vdd FILL
XFILL_9_NOR3X1_33 gnd vdd FILL
XFILL_21_DFFSR_176 gnd vdd FILL
XFILL_2_INVX1_116 gnd vdd FILL
XFILL_9_NOR3X1_44 gnd vdd FILL
XFILL_21_DFFSR_187 gnd vdd FILL
XFILL_21_DFFSR_198 gnd vdd FILL
XFILL_2_INVX1_127 gnd vdd FILL
XFILL_25_DFFSR_120 gnd vdd FILL
XFILL_2_INVX1_138 gnd vdd FILL
XFILL_25_DFFSR_131 gnd vdd FILL
XFILL_2_INVX1_149 gnd vdd FILL
XFILL_25_DFFSR_142 gnd vdd FILL
XFILL_25_DFFSR_153 gnd vdd FILL
XFILL_4_NAND3X1_100 gnd vdd FILL
XFILL_4_NAND3X1_111 gnd vdd FILL
XFILL_25_DFFSR_164 gnd vdd FILL
XFILL_25_DFFSR_175 gnd vdd FILL
XFILL_23_MUX2X1_150 gnd vdd FILL
XFILL_4_NAND3X1_122 gnd vdd FILL
XFILL_23_MUX2X1_161 gnd vdd FILL
XFILL_6_INVX1_104 gnd vdd FILL
XFILL_6_INVX1_115 gnd vdd FILL
XFILL_25_DFFSR_186 gnd vdd FILL
XFILL_23_MUX2X1_172 gnd vdd FILL
XFILL_25_DFFSR_197 gnd vdd FILL
XFILL_6_MUX2X1_110 gnd vdd FILL
XFILL_6_MUX2X1_121 gnd vdd FILL
XFILL_6_INVX1_126 gnd vdd FILL
XFILL_23_MUX2X1_183 gnd vdd FILL
XFILL_29_DFFSR_130 gnd vdd FILL
XFILL_6_INVX1_137 gnd vdd FILL
XFILL_23_MUX2X1_194 gnd vdd FILL
XFILL_6_MUX2X1_132 gnd vdd FILL
XFILL_6_MUX2X1_143 gnd vdd FILL
XFILL_6_INVX1_148 gnd vdd FILL
XFILL_6_INVX1_159 gnd vdd FILL
XFILL_29_DFFSR_141 gnd vdd FILL
XFILL_29_DFFSR_152 gnd vdd FILL
XFILL_6_MUX2X1_154 gnd vdd FILL
XFILL_6_MUX2X1_165 gnd vdd FILL
XFILL_29_DFFSR_163 gnd vdd FILL
XFILL_29_DFFSR_174 gnd vdd FILL
XFILL_6_MUX2X1_176 gnd vdd FILL
XFILL_21_NOR3X1_10 gnd vdd FILL
XFILL_6_MUX2X1_187 gnd vdd FILL
XFILL_29_DFFSR_185 gnd vdd FILL
XFILL_21_NOR3X1_21 gnd vdd FILL
XFILL_21_NOR3X1_32 gnd vdd FILL
XFILL_29_DFFSR_196 gnd vdd FILL
XFILL_21_NOR3X1_43 gnd vdd FILL
XFILL_71_DFFSR_210 gnd vdd FILL
XFILL_54_5_1 gnd vdd FILL
XFILL_71_DFFSR_221 gnd vdd FILL
XFILL_71_DFFSR_232 gnd vdd FILL
XFILL_53_0_0 gnd vdd FILL
XFILL_71_DFFSR_243 gnd vdd FILL
XFILL_71_DFFSR_254 gnd vdd FILL
XFILL_71_DFFSR_265 gnd vdd FILL
XFILL_25_NOR3X1_20 gnd vdd FILL
XFILL_25_NOR3X1_31 gnd vdd FILL
XFILL_25_NOR3X1_42 gnd vdd FILL
XFILL_75_DFFSR_220 gnd vdd FILL
XFILL_75_DFFSR_231 gnd vdd FILL
XFILL_75_DFFSR_242 gnd vdd FILL
XFILL_10_BUFX4_7 gnd vdd FILL
XFILL_75_DFFSR_253 gnd vdd FILL
XFILL_75_DFFSR_264 gnd vdd FILL
XFILL_75_DFFSR_275 gnd vdd FILL
XFILL_30_CLKBUF1_5 gnd vdd FILL
XFILL_29_NOR3X1_30 gnd vdd FILL
XFILL_29_NOR3X1_41 gnd vdd FILL
XFILL_29_NOR3X1_52 gnd vdd FILL
XFILL_79_DFFSR_230 gnd vdd FILL
XFILL_8_OAI22X1_9 gnd vdd FILL
XFILL_79_DFFSR_241 gnd vdd FILL
XFILL_79_DFFSR_252 gnd vdd FILL
XFILL_79_DFFSR_263 gnd vdd FILL
XFILL_79_DFFSR_274 gnd vdd FILL
XFILL_34_CLKBUF1_4 gnd vdd FILL
XFILL_9_NAND3X1_13 gnd vdd FILL
XFILL_9_NAND3X1_24 gnd vdd FILL
XFILL_9_NAND3X1_35 gnd vdd FILL
XFILL_9_NAND3X1_46 gnd vdd FILL
XFILL_9_NAND3X1_57 gnd vdd FILL
XFILL_9_NAND3X1_68 gnd vdd FILL
XFILL_15_BUFX4_15 gnd vdd FILL
XFILL_9_NAND3X1_79 gnd vdd FILL
XFILL_0_NOR3X1_1 gnd vdd FILL
XFILL_15_BUFX4_26 gnd vdd FILL
XFILL_15_BUFX4_37 gnd vdd FILL
XFILL_57_DFFSR_209 gnd vdd FILL
XFILL_15_BUFX4_48 gnd vdd FILL
XFILL_15_BUFX4_59 gnd vdd FILL
XFILL_84_DFFSR_109 gnd vdd FILL
XFILL_2_NAND2X1_15 gnd vdd FILL
XFILL_2_NAND2X1_26 gnd vdd FILL
XFILL_33_DFFSR_1 gnd vdd FILL
XFILL_45_5_1 gnd vdd FILL
XFILL_2_NAND2X1_37 gnd vdd FILL
XFILL_2_NAND2X1_48 gnd vdd FILL
XFILL_44_0_0 gnd vdd FILL
XFILL_2_NAND2X1_59 gnd vdd FILL
XFILL_12_MUX2X1_190 gnd vdd FILL
XFILL_42_DFFSR_220 gnd vdd FILL
XFILL_42_DFFSR_231 gnd vdd FILL
XFILL_42_DFFSR_242 gnd vdd FILL
XFILL_42_DFFSR_253 gnd vdd FILL
XFILL_42_DFFSR_264 gnd vdd FILL
XFILL_42_DFFSR_275 gnd vdd FILL
XFILL_1_NOR2X1_90 gnd vdd FILL
XFILL_28_CLKBUF1_14 gnd vdd FILL
XFILL_28_CLKBUF1_25 gnd vdd FILL
XFILL_55_DFFSR_5 gnd vdd FILL
XFILL_28_CLKBUF1_36 gnd vdd FILL
XFILL_46_DFFSR_230 gnd vdd FILL
XFILL_46_DFFSR_241 gnd vdd FILL
XFILL_7_BUFX4_14 gnd vdd FILL
XFILL_7_BUFX4_25 gnd vdd FILL
XFILL_46_DFFSR_252 gnd vdd FILL
XFILL_7_BUFX4_36 gnd vdd FILL
XFILL_7_BUFX4_47 gnd vdd FILL
XFILL_46_DFFSR_263 gnd vdd FILL
XFILL_46_DFFSR_274 gnd vdd FILL
XFILL_7_BUFX4_58 gnd vdd FILL
XFILL_7_BUFX4_69 gnd vdd FILL
XFILL_6_AOI21X1_15 gnd vdd FILL
XFILL_73_DFFSR_130 gnd vdd FILL
XFILL_6_AOI21X1_26 gnd vdd FILL
XFILL_6_AOI21X1_37 gnd vdd FILL
XFILL_73_DFFSR_141 gnd vdd FILL
XFILL_73_DFFSR_152 gnd vdd FILL
XFILL_73_DFFSR_163 gnd vdd FILL
XFILL_6_AOI21X1_48 gnd vdd FILL
XFILL_6_AOI21X1_59 gnd vdd FILL
XFILL_73_DFFSR_174 gnd vdd FILL
XFILL_16_OAI22X1_17 gnd vdd FILL
XFILL_6_1 gnd vdd FILL
XFILL_16_OAI22X1_28 gnd vdd FILL
XFILL_73_DFFSR_185 gnd vdd FILL
XFILL_16_OAI22X1_39 gnd vdd FILL
XFILL_73_DFFSR_196 gnd vdd FILL
XFILL_9_NOR2X1_103 gnd vdd FILL
XFILL_24_DFFSR_209 gnd vdd FILL
XFILL_9_NOR2X1_114 gnd vdd FILL
XFILL_9_NOR2X1_125 gnd vdd FILL
XFILL_62_3 gnd vdd FILL
XFILL_77_DFFSR_140 gnd vdd FILL
XFILL_77_DFFSR_151 gnd vdd FILL
XFILL_9_NOR2X1_136 gnd vdd FILL
XFILL_77_DFFSR_162 gnd vdd FILL
XFILL_9_NOR2X1_147 gnd vdd FILL
XFILL_0_CLKBUF1_18 gnd vdd FILL
XFILL_9_NOR2X1_158 gnd vdd FILL
XFILL_77_DFFSR_173 gnd vdd FILL
XFILL_77_DFFSR_184 gnd vdd FILL
XFILL_0_CLKBUF1_29 gnd vdd FILL
XFILL_9_NOR2X1_169 gnd vdd FILL
XFILL_51_DFFSR_109 gnd vdd FILL
XFILL_77_DFFSR_9 gnd vdd FILL
XFILL_15_NAND3X1_60 gnd vdd FILL
XFILL_77_DFFSR_195 gnd vdd FILL
XFILL_15_NAND3X1_71 gnd vdd FILL
XFILL_28_DFFSR_208 gnd vdd FILL
XFILL_14_AND2X2_2 gnd vdd FILL
XFILL_28_DFFSR_219 gnd vdd FILL
XFILL_15_NAND3X1_82 gnd vdd FILL
XFILL_15_NAND3X1_93 gnd vdd FILL
XFILL_36_5_1 gnd vdd FILL
XFILL_35_0_0 gnd vdd FILL
XFILL_1_NAND2X1_1 gnd vdd FILL
XFILL_55_DFFSR_108 gnd vdd FILL
XFILL_55_DFFSR_119 gnd vdd FILL
XFILL_11_BUFX4_30 gnd vdd FILL
XFILL_11_BUFX4_41 gnd vdd FILL
XFILL_59_DFFSR_107 gnd vdd FILL
XFILL_9_MUX2X1_109 gnd vdd FILL
XFILL_11_BUFX4_52 gnd vdd FILL
XFILL_59_DFFSR_118 gnd vdd FILL
XFILL_11_BUFX4_63 gnd vdd FILL
XFILL_59_DFFSR_129 gnd vdd FILL
XFILL_11_BUFX4_74 gnd vdd FILL
XFILL_11_BUFX4_85 gnd vdd FILL
XFILL_11_BUFX4_96 gnd vdd FILL
XFILL_6_OAI22X1_12 gnd vdd FILL
XFILL_6_OAI22X1_23 gnd vdd FILL
XFILL_6_OAI22X1_34 gnd vdd FILL
XDFFSR_11 INVX1_31/A DFFSR_8/CLK DFFSR_8/R vdd DFFSR_11/D gnd vdd DFFSR
XFILL_6_OAI22X1_45 gnd vdd FILL
XFILL_60_DFFSR_19 gnd vdd FILL
XDFFSR_22 DFFSR_22/Q DFFSR_88/CLK DFFSR_87/R vdd DFFSR_22/D gnd vdd DFFSR
XDFFSR_33 INVX1_26/A DFFSR_79/CLK DFFSR_79/R vdd DFFSR_33/D gnd vdd DFFSR
XDFFSR_44 INVX1_20/A CLKBUF1_5/Y DFFSR_49/R vdd MUX2X1_7/Y gnd vdd DFFSR
XDFFSR_55 INVX1_4/A DFFSR_55/CLK DFFSR_55/R vdd DFFSR_55/D gnd vdd DFFSR
XDFFSR_66 DFFSR_66/Q DFFSR_76/CLK DFFSR_97/R vdd DFFSR_66/D gnd vdd DFFSR
XFILL_13_DFFSR_230 gnd vdd FILL
XFILL_13_DFFSR_241 gnd vdd FILL
XDFFSR_77 DFFSR_77/Q CLKBUF1_8/Y DFFSR_82/R vdd DFFSR_77/D gnd vdd DFFSR
XDFFSR_88 DFFSR_88/Q DFFSR_88/CLK DFFSR_91/R vdd DFFSR_88/D gnd vdd DFFSR
XFILL_13_DFFSR_252 gnd vdd FILL
XDFFSR_99 DFFSR_99/Q DFFSR_99/CLK DFFSR_99/R vdd DFFSR_99/D gnd vdd DFFSR
XFILL_13_DFFSR_263 gnd vdd FILL
XFILL_13_DFFSR_274 gnd vdd FILL
XFILL_10_MUX2X1_19 gnd vdd FILL
XFILL_3_NOR2X1_203 gnd vdd FILL
XFILL_40_DFFSR_130 gnd vdd FILL
XFILL_1_AOI21X1_6 gnd vdd FILL
XFILL_17_DFFSR_240 gnd vdd FILL
XFILL_40_DFFSR_141 gnd vdd FILL
XFILL_5_INVX1_20 gnd vdd FILL
XFILL_40_DFFSR_152 gnd vdd FILL
XFILL_5_INVX1_31 gnd vdd FILL
XFILL_5_NAND3X1_101 gnd vdd FILL
XFILL_9_NAND2X1_90 gnd vdd FILL
XFILL_14_BUFX4_8 gnd vdd FILL
XCLKBUF1_20 BUFX4_95/Y gnd DFFSR_56/CLK vdd CLKBUF1
XFILL_17_DFFSR_251 gnd vdd FILL
XFILL_40_DFFSR_163 gnd vdd FILL
XFILL_5_NAND3X1_112 gnd vdd FILL
XFILL_17_DFFSR_262 gnd vdd FILL
XCLKBUF1_31 BUFX4_73/Y gnd CLKBUF1_31/Y vdd CLKBUF1
XFILL_5_INVX1_42 gnd vdd FILL
XFILL_5_NAND3X1_123 gnd vdd FILL
XFILL_6_AND2X2_1 gnd vdd FILL
XFILL_40_DFFSR_174 gnd vdd FILL
XFILL_5_INVX1_53 gnd vdd FILL
XCLKBUF1_42 BUFX4_73/Y gnd DFFSR_64/CLK vdd CLKBUF1
XFILL_17_DFFSR_273 gnd vdd FILL
XFILL_5_INVX1_64 gnd vdd FILL
XFILL_14_MUX2X1_18 gnd vdd FILL
XFILL_40_DFFSR_185 gnd vdd FILL
XFILL_5_INVX1_75 gnd vdd FILL
XFILL_17_CLKBUF1_10 gnd vdd FILL
XFILL_40_DFFSR_196 gnd vdd FILL
XFILL_17_CLKBUF1_21 gnd vdd FILL
XFILL_5_INVX1_86 gnd vdd FILL
XFILL_14_MUX2X1_29 gnd vdd FILL
XFILL_17_CLKBUF1_32 gnd vdd FILL
XFILL_5_INVX1_97 gnd vdd FILL
XFILL_5_AOI21X1_5 gnd vdd FILL
XFILL_44_DFFSR_140 gnd vdd FILL
XFILL_44_DFFSR_151 gnd vdd FILL
XFILL_44_DFFSR_162 gnd vdd FILL
XFILL_44_DFFSR_173 gnd vdd FILL
XFILL_12_MUX2X1_7 gnd vdd FILL
XFILL_12_AOI21X1_40 gnd vdd FILL
XFILL_44_DFFSR_184 gnd vdd FILL
XFILL_12_AOI21X1_51 gnd vdd FILL
XFILL_2_5_1 gnd vdd FILL
XFILL_18_MUX2X1_17 gnd vdd FILL
XFILL_27_5_1 gnd vdd FILL
XFILL_44_DFFSR_195 gnd vdd FILL
XFILL_12_AOI21X1_62 gnd vdd FILL
XFILL_18_MUX2X1_28 gnd vdd FILL
XFILL_12_AOI21X1_73 gnd vdd FILL
XFILL_26_0_0 gnd vdd FILL
XFILL_18_MUX2X1_39 gnd vdd FILL
XFILL_1_0_0 gnd vdd FILL
XFILL_9_AOI21X1_4 gnd vdd FILL
XFILL_48_DFFSR_150 gnd vdd FILL
XFILL_3_BUFX4_40 gnd vdd FILL
XFILL_10_AOI22X1_2 gnd vdd FILL
XFILL_48_DFFSR_161 gnd vdd FILL
XFILL_3_BUFX4_51 gnd vdd FILL
XFILL_48_DFFSR_172 gnd vdd FILL
XFILL_3_BUFX4_62 gnd vdd FILL
XFILL_3_BUFX4_73 gnd vdd FILL
XFILL_48_DFFSR_183 gnd vdd FILL
XFILL_3_BUFX4_84 gnd vdd FILL
XFILL_22_DFFSR_108 gnd vdd FILL
XFILL_48_DFFSR_194 gnd vdd FILL
XFILL_3_BUFX4_95 gnd vdd FILL
XFILL_22_DFFSR_119 gnd vdd FILL
XFILL_10_BUFX2_4 gnd vdd FILL
XFILL_14_AOI22X1_1 gnd vdd FILL
XFILL_10_4_1 gnd vdd FILL
XFILL_26_DFFSR_107 gnd vdd FILL
XFILL_26_DFFSR_118 gnd vdd FILL
XFILL_21_MUX2X1_5 gnd vdd FILL
XFILL_26_DFFSR_129 gnd vdd FILL
XINVX1_105 INVX1_105/A gnd MUX2X1_92/A vdd INVX1
XFILL_0_NAND3X1_130 gnd vdd FILL
XFILL_37_DFFSR_2 gnd vdd FILL
XINVX1_116 DFFSR_24/Q gnd NOR3X1_26/A vdd INVX1
XINVX1_127 OAI22X1_3/D gnd INVX1_127/Y vdd INVX1
XFILL_5_NOR2X1_8 gnd vdd FILL
XINVX1_138 AND2X2_2/A gnd INVX1_138/Y vdd INVX1
XFILL_29_DFFSR_20 gnd vdd FILL
XFILL_15_MUX2X1_101 gnd vdd FILL
XFILL_29_DFFSR_31 gnd vdd FILL
XINVX1_149 INVX1_149/A gnd INVX1_149/Y vdd INVX1
XFILL_15_MUX2X1_112 gnd vdd FILL
XFILL_15_MUX2X1_123 gnd vdd FILL
XFILL_29_DFFSR_42 gnd vdd FILL
XFILL_29_DFFSR_53 gnd vdd FILL
XFILL_29_DFFSR_64 gnd vdd FILL
XFILL_15_MUX2X1_134 gnd vdd FILL
XFILL_15_MUX2X1_145 gnd vdd FILL
XFILL_29_DFFSR_75 gnd vdd FILL
XFILL_15_MUX2X1_156 gnd vdd FILL
XFILL_29_DFFSR_86 gnd vdd FILL
XFILL_9_1_0 gnd vdd FILL
XFILL_15_MUX2X1_167 gnd vdd FILL
XFILL_22_NOR3X1_19 gnd vdd FILL
XFILL_15_MUX2X1_178 gnd vdd FILL
XFILL_29_DFFSR_97 gnd vdd FILL
XFILL_15_MUX2X1_189 gnd vdd FILL
XFILL_69_DFFSR_30 gnd vdd FILL
XFILL_72_DFFSR_208 gnd vdd FILL
XFILL_69_DFFSR_41 gnd vdd FILL
XFILL_72_DFFSR_219 gnd vdd FILL
XFILL_4_MUX2X1_6 gnd vdd FILL
XFILL_69_DFFSR_52 gnd vdd FILL
XFILL_69_DFFSR_63 gnd vdd FILL
XFILL_69_DFFSR_74 gnd vdd FILL
XFILL_21_DFFSR_8 gnd vdd FILL
XFILL_69_DFFSR_85 gnd vdd FILL
XFILL_26_NOR3X1_18 gnd vdd FILL
XFILL_69_DFFSR_96 gnd vdd FILL
XFILL_26_NOR3X1_29 gnd vdd FILL
XFILL_76_DFFSR_207 gnd vdd FILL
XFILL_59_DFFSR_6 gnd vdd FILL
XFILL_76_DFFSR_218 gnd vdd FILL
XFILL_11_DFFSR_140 gnd vdd FILL
XFILL_18_5_1 gnd vdd FILL
XFILL_76_DFFSR_229 gnd vdd FILL
XFILL_11_DFFSR_151 gnd vdd FILL
XFILL_11_DFFSR_162 gnd vdd FILL
XFILL_38_DFFSR_40 gnd vdd FILL
XFILL_11_DFFSR_173 gnd vdd FILL
XFILL_17_0_0 gnd vdd FILL
XFILL_38_DFFSR_51 gnd vdd FILL
XFILL_0_CLKBUF1_5 gnd vdd FILL
XFILL_11_DFFSR_184 gnd vdd FILL
XFILL_38_DFFSR_62 gnd vdd FILL
XFILL_11_DFFSR_195 gnd vdd FILL
XFILL_38_DFFSR_73 gnd vdd FILL
XFILL_38_DFFSR_84 gnd vdd FILL
XFILL_38_DFFSR_95 gnd vdd FILL
XFILL_60_3_1 gnd vdd FILL
XFILL_15_DFFSR_150 gnd vdd FILL
XFILL_27_6 gnd vdd FILL
XFILL_15_DFFSR_161 gnd vdd FILL
XFILL_15_DFFSR_172 gnd vdd FILL
XFILL_4_CLKBUF1_4 gnd vdd FILL
XFILL_78_DFFSR_50 gnd vdd FILL
XFILL_15_DFFSR_183 gnd vdd FILL
XFILL_78_DFFSR_61 gnd vdd FILL
XFILL_15_DFFSR_194 gnd vdd FILL
XFILL_22_MUX2X1_180 gnd vdd FILL
XFILL_78_DFFSR_72 gnd vdd FILL
XFILL_78_DFFSR_83 gnd vdd FILL
XFILL_22_MUX2X1_191 gnd vdd FILL
XFILL_5_MUX2X1_140 gnd vdd FILL
XFILL_78_DFFSR_94 gnd vdd FILL
XFILL_5_MUX2X1_151 gnd vdd FILL
XFILL_19_DFFSR_160 gnd vdd FILL
XFILL_5_MUX2X1_162 gnd vdd FILL
XFILL_8_CLKBUF1_3 gnd vdd FILL
XFILL_5_MUX2X1_173 gnd vdd FILL
XFILL_19_DFFSR_171 gnd vdd FILL
XFILL_5_MUX2X1_184 gnd vdd FILL
XFILL_19_DFFSR_182 gnd vdd FILL
XFILL_19_DFFSR_193 gnd vdd FILL
XFILL_1_INVX1_90 gnd vdd FILL
XFILL_18_NOR3X1_2 gnd vdd FILL
XFILL_11_NOR3X1_40 gnd vdd FILL
XFILL_1_BUFX2_10 gnd vdd FILL
XFILL_11_NOR3X1_51 gnd vdd FILL
XFILL_47_DFFSR_60 gnd vdd FILL
XFILL_47_DFFSR_71 gnd vdd FILL
XFILL_61_DFFSR_240 gnd vdd FILL
XFILL_47_DFFSR_82 gnd vdd FILL
XFILL_47_DFFSR_93 gnd vdd FILL
XFILL_61_DFFSR_251 gnd vdd FILL
XFILL_61_DFFSR_262 gnd vdd FILL
XFILL_61_DFFSR_273 gnd vdd FILL
XFILL_15_NOR3X1_50 gnd vdd FILL
XFILL_87_DFFSR_70 gnd vdd FILL
XFILL_87_DFFSR_81 gnd vdd FILL
XFILL_65_DFFSR_250 gnd vdd FILL
XFILL_87_DFFSR_92 gnd vdd FILL
XFILL_65_DFFSR_261 gnd vdd FILL
XFILL_65_DFFSR_272 gnd vdd FILL
XFILL_16_DFFSR_70 gnd vdd FILL
XFILL_20_CLKBUF1_2 gnd vdd FILL
XFILL_11_NAND2X1_17 gnd vdd FILL
XFILL_16_DFFSR_81 gnd vdd FILL
XFILL_11_NAND2X1_28 gnd vdd FILL
XFILL_16_DFFSR_92 gnd vdd FILL
XFILL_11_NAND2X1_39 gnd vdd FILL
XFILL_1_OAI21X1_9 gnd vdd FILL
XFILL_69_DFFSR_260 gnd vdd FILL
XFILL_24_CLKBUF1_1 gnd vdd FILL
XFILL_69_DFFSR_271 gnd vdd FILL
XFILL_56_DFFSR_80 gnd vdd FILL
XFILL_56_DFFSR_91 gnd vdd FILL
XFILL_2_NOR2X1_11 gnd vdd FILL
XFILL_43_DFFSR_207 gnd vdd FILL
XFILL_8_NAND3X1_10 gnd vdd FILL
XFILL_2_NOR2X1_22 gnd vdd FILL
XFILL_8_NAND3X1_21 gnd vdd FILL
XFILL_2_NOR2X1_33 gnd vdd FILL
XFILL_43_DFFSR_218 gnd vdd FILL
XFILL_5_OAI21X1_8 gnd vdd FILL
XFILL_43_DFFSR_229 gnd vdd FILL
XFILL_2_NOR2X1_44 gnd vdd FILL
XFILL_8_NAND3X1_32 gnd vdd FILL
XFILL_1_NOR2X1_1 gnd vdd FILL
XFILL_2_NOR2X1_55 gnd vdd FILL
XFILL_8_NAND3X1_43 gnd vdd FILL
XFILL_2_NOR2X1_66 gnd vdd FILL
XFILL_8_NAND3X1_54 gnd vdd FILL
XFILL_8_NAND3X1_65 gnd vdd FILL
XFILL_2_NOR2X1_77 gnd vdd FILL
XFILL_51_3_1 gnd vdd FILL
XFILL_8_NAND3X1_76 gnd vdd FILL
XFILL_2_NOR2X1_88 gnd vdd FILL
XFILL_70_DFFSR_107 gnd vdd FILL
XFILL_8_NAND3X1_87 gnd vdd FILL
XFILL_2_NOR2X1_99 gnd vdd FILL
XFILL_6_NOR2X1_10 gnd vdd FILL
XFILL_47_DFFSR_206 gnd vdd FILL
XFILL_70_DFFSR_118 gnd vdd FILL
XFILL_6_NOR2X1_21 gnd vdd FILL
XFILL_8_NAND3X1_98 gnd vdd FILL
XFILL_47_DFFSR_217 gnd vdd FILL
XFILL_6_NOR2X1_32 gnd vdd FILL
XFILL_9_OAI21X1_7 gnd vdd FILL
XFILL_47_DFFSR_228 gnd vdd FILL
XFILL_70_DFFSR_129 gnd vdd FILL
XFILL_6_NOR2X1_43 gnd vdd FILL
XFILL_47_DFFSR_239 gnd vdd FILL
XFILL_25_DFFSR_90 gnd vdd FILL
XFILL_6_NOR2X1_54 gnd vdd FILL
XFILL_10_OAI22X1_5 gnd vdd FILL
XFILL_6_NOR2X1_65 gnd vdd FILL
XFILL_6_NOR2X1_76 gnd vdd FILL
XFILL_6_NOR2X1_87 gnd vdd FILL
XFILL_74_DFFSR_106 gnd vdd FILL
XFILL_6_NOR2X1_98 gnd vdd FILL
XFILL_74_DFFSR_117 gnd vdd FILL
XFILL_74_DFFSR_128 gnd vdd FILL
XFILL_74_DFFSR_139 gnd vdd FILL
XFILL_14_OAI22X1_4 gnd vdd FILL
XFILL_15_AOI21X1_17 gnd vdd FILL
XFILL_15_AOI21X1_28 gnd vdd FILL
XFILL_1_NAND2X1_12 gnd vdd FILL
XFILL_1_NAND2X1_23 gnd vdd FILL
XFILL_6_DFFSR_1 gnd vdd FILL
XFILL_15_AOI21X1_39 gnd vdd FILL
XFILL_1_NAND2X1_34 gnd vdd FILL
XFILL_15_NAND3X1_130 gnd vdd FILL
XFILL_1_NAND2X1_45 gnd vdd FILL
XFILL_78_DFFSR_105 gnd vdd FILL
XFILL_78_DFFSR_116 gnd vdd FILL
XFILL_1_NAND2X1_56 gnd vdd FILL
XFILL_78_DFFSR_127 gnd vdd FILL
XFILL_12_BUFX4_19 gnd vdd FILL
XFILL_1_NAND2X1_67 gnd vdd FILL
XFILL_1_NAND2X1_78 gnd vdd FILL
XFILL_78_DFFSR_138 gnd vdd FILL
XFILL_1_NAND2X1_89 gnd vdd FILL
XFILL_78_DFFSR_149 gnd vdd FILL
XFILL_18_OAI22X1_3 gnd vdd FILL
XFILL_8_DFFSR_80 gnd vdd FILL
XFILL_8_DFFSR_91 gnd vdd FILL
XFILL_1_BUFX2_7 gnd vdd FILL
XFILL_59_4_1 gnd vdd FILL
XFILL_6_NAND3X1_102 gnd vdd FILL
XFILL_6_NAND3X1_113 gnd vdd FILL
XFILL_32_DFFSR_250 gnd vdd FILL
XFILL_6_NAND3X1_124 gnd vdd FILL
XFILL_32_DFFSR_261 gnd vdd FILL
XFILL_32_DFFSR_272 gnd vdd FILL
XFILL_27_CLKBUF1_11 gnd vdd FILL
XFILL_27_CLKBUF1_22 gnd vdd FILL
XFILL_60_DFFSR_6 gnd vdd FILL
XFILL_27_CLKBUF1_33 gnd vdd FILL
XFILL_1_AOI22X1_10 gnd vdd FILL
XFILL_36_DFFSR_260 gnd vdd FILL
XFILL_36_DFFSR_271 gnd vdd FILL
XFILL_12_OR2X2_1 gnd vdd FILL
XFILL_6_NAND2X1_9 gnd vdd FILL
XFILL_10_DFFSR_207 gnd vdd FILL
XFILL_2_MUX2X1_40 gnd vdd FILL
XFILL_2_MUX2X1_51 gnd vdd FILL
XFILL_5_AOI21X1_12 gnd vdd FILL
XFILL_10_DFFSR_218 gnd vdd FILL
XFILL_2_MUX2X1_62 gnd vdd FILL
XFILL_10_DFFSR_229 gnd vdd FILL
XFILL_5_AOI21X1_23 gnd vdd FILL
XFILL_5_AOI21X1_34 gnd vdd FILL
XFILL_2_MUX2X1_73 gnd vdd FILL
XFILL_42_3_1 gnd vdd FILL
XFILL_5_AOI21X1_45 gnd vdd FILL
XFILL_2_MUX2X1_84 gnd vdd FILL
XFILL_63_DFFSR_160 gnd vdd FILL
XFILL_2_MUX2X1_95 gnd vdd FILL
XFILL_15_OAI22X1_14 gnd vdd FILL
XFILL_5_AOI21X1_56 gnd vdd FILL
XFILL_63_DFFSR_171 gnd vdd FILL
XFILL_5_AOI21X1_67 gnd vdd FILL
XFILL_15_OAI22X1_25 gnd vdd FILL
XFILL_63_DFFSR_182 gnd vdd FILL
XFILL_5_AOI21X1_78 gnd vdd FILL
XFILL_63_DFFSR_193 gnd vdd FILL
XFILL_15_OAI22X1_36 gnd vdd FILL
XFILL_14_DFFSR_206 gnd vdd FILL
XFILL_15_OAI22X1_47 gnd vdd FILL
XFILL_11_NAND3X1_6 gnd vdd FILL
XFILL_8_NOR2X1_100 gnd vdd FILL
XFILL_14_DFFSR_217 gnd vdd FILL
XFILL_8_NOR2X1_111 gnd vdd FILL
XFILL_6_MUX2X1_50 gnd vdd FILL
XFILL_14_DFFSR_228 gnd vdd FILL
XFILL_6_MUX2X1_61 gnd vdd FILL
XFILL_8_NOR2X1_122 gnd vdd FILL
XFILL_8_NOR2X1_133 gnd vdd FILL
XFILL_14_DFFSR_239 gnd vdd FILL
XFILL_6_MUX2X1_72 gnd vdd FILL
XFILL_6_MUX2X1_83 gnd vdd FILL
XFILL_0_BUFX4_1 gnd vdd FILL
XFILL_6_MUX2X1_94 gnd vdd FILL
XFILL_8_NOR2X1_144 gnd vdd FILL
XFILL_25_DFFSR_9 gnd vdd FILL
XFILL_67_DFFSR_170 gnd vdd FILL
XFILL_8_NOR2X1_155 gnd vdd FILL
XFILL_4_BUFX4_18 gnd vdd FILL
XFILL_8_NOR2X1_166 gnd vdd FILL
XFILL_67_DFFSR_181 gnd vdd FILL
XFILL_4_BUFX4_29 gnd vdd FILL
XFILL_8_NOR2X1_177 gnd vdd FILL
XFILL_67_DFFSR_192 gnd vdd FILL
XFILL_41_DFFSR_106 gnd vdd FILL
XFILL_8_NOR2X1_188 gnd vdd FILL
XFILL_18_DFFSR_205 gnd vdd FILL
XFILL_41_DFFSR_117 gnd vdd FILL
XFILL_15_NAND3X1_5 gnd vdd FILL
XFILL_8_NOR2X1_199 gnd vdd FILL
XFILL_18_DFFSR_216 gnd vdd FILL
XFILL_18_DFFSR_227 gnd vdd FILL
XFILL_41_DFFSR_128 gnd vdd FILL
XFILL_14_NAND3X1_90 gnd vdd FILL
XFILL_18_DFFSR_238 gnd vdd FILL
XFILL_41_DFFSR_139 gnd vdd FILL
XFILL_18_DFFSR_249 gnd vdd FILL
XFILL_1_NAND3X1_120 gnd vdd FILL
XFILL_1_NAND3X1_131 gnd vdd FILL
XFILL_45_DFFSR_105 gnd vdd FILL
XFILL_45_DFFSR_116 gnd vdd FILL
XFILL_45_DFFSR_127 gnd vdd FILL
XFILL_45_DFFSR_138 gnd vdd FILL
XFILL_45_DFFSR_149 gnd vdd FILL
XFILL_49_DFFSR_104 gnd vdd FILL
XFILL_8_MUX2X1_106 gnd vdd FILL
XFILL_8_MUX2X1_117 gnd vdd FILL
XFILL_49_DFFSR_115 gnd vdd FILL
XFILL_49_DFFSR_126 gnd vdd FILL
XFILL_8_MUX2X1_128 gnd vdd FILL
XFILL_49_DFFSR_137 gnd vdd FILL
XFILL_8_MUX2X1_139 gnd vdd FILL
XFILL_49_DFFSR_148 gnd vdd FILL
XFILL_11_AND2X2_6 gnd vdd FILL
XFILL_22_MUX2X1_70 gnd vdd FILL
XFILL_5_OAI22X1_20 gnd vdd FILL
XFILL_49_DFFSR_159 gnd vdd FILL
XFILL_22_MUX2X1_81 gnd vdd FILL
XFILL_5_OAI22X1_31 gnd vdd FILL
XFILL_5_OAI22X1_42 gnd vdd FILL
XFILL_22_MUX2X1_92 gnd vdd FILL
XFILL_9_OAI21X1_11 gnd vdd FILL
XFILL_9_OAI21X1_22 gnd vdd FILL
XFILL_9_OAI21X1_33 gnd vdd FILL
XFILL_9_OAI21X1_44 gnd vdd FILL
XFILL_0_INVX4_1 gnd vdd FILL
XFILL_32_4 gnd vdd FILL
XFILL_33_3_1 gnd vdd FILL
XFILL_2_NOR2X1_200 gnd vdd FILL
XFILL_25_3 gnd vdd FILL
XFILL_19_AOI22X1_9 gnd vdd FILL
XFILL_30_DFFSR_160 gnd vdd FILL
XFILL_18_2 gnd vdd FILL
XFILL_30_DFFSR_171 gnd vdd FILL
XFILL_30_DFFSR_182 gnd vdd FILL
XFILL_30_DFFSR_193 gnd vdd FILL
XFILL_39_DFFSR_18 gnd vdd FILL
XFILL_39_DFFSR_29 gnd vdd FILL
XFILL_16_CLKBUF1_40 gnd vdd FILL
XFILL_34_DFFSR_170 gnd vdd FILL
XFILL_34_DFFSR_181 gnd vdd FILL
XFILL_79_DFFSR_17 gnd vdd FILL
XFILL_34_DFFSR_192 gnd vdd FILL
XFILL_11_AOI21X1_70 gnd vdd FILL
XFILL_79_DFFSR_28 gnd vdd FILL
XFILL_11_AOI21X1_81 gnd vdd FILL
XFILL_79_DFFSR_39 gnd vdd FILL
XFILL_2_INVX1_13 gnd vdd FILL
XFILL_38_DFFSR_180 gnd vdd FILL
XFILL_2_INVX1_24 gnd vdd FILL
XFILL_2_INVX1_35 gnd vdd FILL
XFILL_38_DFFSR_191 gnd vdd FILL
XFILL_12_DFFSR_105 gnd vdd FILL
XFILL_2_INVX1_46 gnd vdd FILL
XFILL_3_AND2X2_5 gnd vdd FILL
XFILL_12_DFFSR_116 gnd vdd FILL
XFILL_2_INVX1_57 gnd vdd FILL
XFILL_12_DFFSR_127 gnd vdd FILL
XFILL_2_INVX1_68 gnd vdd FILL
XFILL_12_DFFSR_138 gnd vdd FILL
XFILL_2_INVX1_79 gnd vdd FILL
XFILL_12_DFFSR_149 gnd vdd FILL
XFILL_48_DFFSR_16 gnd vdd FILL
XFILL_48_DFFSR_27 gnd vdd FILL
XFILL_48_DFFSR_38 gnd vdd FILL
XFILL_48_DFFSR_49 gnd vdd FILL
XFILL_80_DFFSR_260 gnd vdd FILL
XFILL_16_DFFSR_104 gnd vdd FILL
XFILL_80_DFFSR_271 gnd vdd FILL
XFILL_16_DFFSR_115 gnd vdd FILL
XFILL_16_DFFSR_126 gnd vdd FILL
XFILL_16_DFFSR_137 gnd vdd FILL
XFILL_0_BUFX4_11 gnd vdd FILL
XFILL_16_DFFSR_148 gnd vdd FILL
XFILL_42_DFFSR_3 gnd vdd FILL
XFILL_0_BUFX4_22 gnd vdd FILL
XFILL_16_DFFSR_159 gnd vdd FILL
XFILL_0_BUFX4_33 gnd vdd FILL
XFILL_0_BUFX4_44 gnd vdd FILL
XFILL_17_DFFSR_15 gnd vdd FILL
XFILL_84_DFFSR_270 gnd vdd FILL
XFILL_0_BUFX4_55 gnd vdd FILL
XFILL_17_DFFSR_26 gnd vdd FILL
XFILL_0_BUFX4_66 gnd vdd FILL
XFILL_17_DFFSR_37 gnd vdd FILL
XFILL_0_BUFX4_77 gnd vdd FILL
XFILL_17_DFFSR_48 gnd vdd FILL
XFILL_14_MUX2X1_120 gnd vdd FILL
XFILL_17_DFFSR_59 gnd vdd FILL
XFILL_0_BUFX4_88 gnd vdd FILL
XFILL_0_BUFX4_99 gnd vdd FILL
XFILL_14_MUX2X1_131 gnd vdd FILL
XFILL_24_3_1 gnd vdd FILL
XFILL_14_MUX2X1_142 gnd vdd FILL
XFILL_14_MUX2X1_153 gnd vdd FILL
XFILL_12_NOR3X1_16 gnd vdd FILL
XFILL_14_MUX2X1_164 gnd vdd FILL
XFILL_57_DFFSR_14 gnd vdd FILL
XFILL_14_MUX2X1_175 gnd vdd FILL
XFILL_5_BUFX2_8 gnd vdd FILL
XFILL_12_NOR3X1_27 gnd vdd FILL
XFILL_57_DFFSR_25 gnd vdd FILL
XFILL_14_MUX2X1_186 gnd vdd FILL
XFILL_12_NOR3X1_38 gnd vdd FILL
XFILL_12_NOR3X1_49 gnd vdd FILL
XFILL_57_DFFSR_36 gnd vdd FILL
XFILL_62_DFFSR_205 gnd vdd FILL
XFILL_57_DFFSR_47 gnd vdd FILL
XFILL_57_DFFSR_58 gnd vdd FILL
XFILL_62_DFFSR_216 gnd vdd FILL
XFILL_62_DFFSR_227 gnd vdd FILL
XFILL_57_DFFSR_69 gnd vdd FILL
XFILL_62_DFFSR_238 gnd vdd FILL
XFILL_62_DFFSR_249 gnd vdd FILL
XFILL_16_NOR3X1_15 gnd vdd FILL
XFILL_16_NOR3X1_26 gnd vdd FILL
XFILL_16_NOR3X1_37 gnd vdd FILL
XFILL_16_NOR3X1_48 gnd vdd FILL
XFILL_66_DFFSR_204 gnd vdd FILL
XFILL_64_DFFSR_7 gnd vdd FILL
XFILL_26_DFFSR_13 gnd vdd FILL
XFILL_66_DFFSR_215 gnd vdd FILL
XFILL_26_DFFSR_24 gnd vdd FILL
XFILL_66_DFFSR_226 gnd vdd FILL
XFILL_26_DFFSR_35 gnd vdd FILL
XFILL_66_DFFSR_237 gnd vdd FILL
XFILL_66_DFFSR_248 gnd vdd FILL
XFILL_26_DFFSR_46 gnd vdd FILL
XFILL_26_DFFSR_57 gnd vdd FILL
XFILL_66_DFFSR_259 gnd vdd FILL
XFILL_26_DFFSR_68 gnd vdd FILL
XFILL_26_DFFSR_79 gnd vdd FILL
XFILL_66_DFFSR_12 gnd vdd FILL
XFILL_66_DFFSR_23 gnd vdd FILL
XFILL_66_DFFSR_34 gnd vdd FILL
XFILL_66_DFFSR_45 gnd vdd FILL
XFILL_66_DFFSR_56 gnd vdd FILL
XFILL_66_DFFSR_67 gnd vdd FILL
XFILL_66_DFFSR_78 gnd vdd FILL
XNAND3X1_11 NAND3X1_11/A NAND3X1_11/B AOI22X1_9/Y gnd NOR3X1_44/A vdd NAND3X1
XFILL_66_DFFSR_89 gnd vdd FILL
XFILL_7_4_1 gnd vdd FILL
XNAND3X1_22 DFFSR_84/Q BUFX4_1/Y NOR2X1_44/Y gnd OAI21X1_30/C vdd NAND3X1
XNAND3X1_33 INVX2_4/A OAI21X1_35/A OAI21X1_48/A gnd NAND3X1_33/Y vdd NAND3X1
XNAND3X1_44 DFFSR_28/Q NAND3X1_7/B NOR2X1_37/Y gnd NAND3X1_46/A vdd NAND3X1
XNAND3X1_55 AOI22X1_6/Y NAND3X1_55/B NOR3X1_7/Y gnd NOR3X1_8/C vdd NAND3X1
XFILL_4_BUFX4_2 gnd vdd FILL
XFILL_9_DFFSR_14 gnd vdd FILL
XNAND3X1_66 OAI22X1_7/D OAI22X1_6/D OAI21X1_49/Y gnd NOR3X1_46/C vdd NAND3X1
XFILL_9_DFFSR_25 gnd vdd FILL
XFILL_9_DFFSR_36 gnd vdd FILL
XFILL_4_MUX2X1_170 gnd vdd FILL
XFILL_7_NAND3X1_103 gnd vdd FILL
XNAND3X1_77 NOR3X1_8/Y NOR3X1_11/Y NOR3X1_3/Y gnd DFFSR_243/D vdd NAND3X1
XFILL_35_DFFSR_11 gnd vdd FILL
XFILL_7_NAND3X1_114 gnd vdd FILL
XFILL_4_MUX2X1_181 gnd vdd FILL
XFILL_29_CLKBUF1_9 gnd vdd FILL
XNAND3X1_88 NOR3X1_24/Y NOR2X1_67/Y NOR3X1_20/Y gnd NOR2X1_74/B vdd NAND3X1
XFILL_35_DFFSR_22 gnd vdd FILL
XFILL_7_NAND3X1_125 gnd vdd FILL
XFILL_4_MUX2X1_192 gnd vdd FILL
XFILL_9_DFFSR_47 gnd vdd FILL
XNAND3X1_99 NOR2X1_26/A BUFX4_60/Y NOR3X1_2/Y gnd NAND3X1_99/Y vdd NAND3X1
XFILL_9_DFFSR_58 gnd vdd FILL
XNOR2X1_11 NOR2X1_11/A NOR2X1_12/B gnd NOR2X1_11/Y vdd NOR2X1
XFILL_35_DFFSR_33 gnd vdd FILL
XFILL_9_DFFSR_69 gnd vdd FILL
XNOR2X1_22 NOR2X1_57/A OR2X2_1/A gnd NOR2X1_22/Y vdd NOR2X1
XFILL_35_DFFSR_44 gnd vdd FILL
XFILL_7_NOR2X1_19 gnd vdd FILL
XFILL_35_DFFSR_55 gnd vdd FILL
XNOR2X1_33 NOR2X1_33/A NOR2X1_33/B gnd NOR2X1_33/Y vdd NOR2X1
XNOR2X1_44 NOR3X1_51/C NOR2X1_44/B gnd NOR2X1_44/Y vdd NOR2X1
XNOR2X1_55 OAI21X1_3/Y OAI21X1_2/Y gnd NOR2X1_55/Y vdd NOR2X1
XFILL_35_DFFSR_66 gnd vdd FILL
XFILL_35_DFFSR_77 gnd vdd FILL
XNOR2X1_66 MUX2X1_9/B NOR2X1_66/B gnd NOR3X1_24/C vdd NOR2X1
XFILL_35_DFFSR_88 gnd vdd FILL
XNOR2X1_77 NOR2X1_77/A NOR2X1_77/B gnd NOR2X1_77/Y vdd NOR2X1
XFILL_35_DFFSR_99 gnd vdd FILL
XFILL_75_DFFSR_10 gnd vdd FILL
XNOR2X1_88 INVX1_74/Y OAI22X1_1/B gnd NOR3X1_32/B vdd NOR2X1
XFILL_75_DFFSR_21 gnd vdd FILL
XNOR2X1_99 NOR2X1_99/A NOR2X1_99/B gnd NOR2X1_99/Y vdd NOR2X1
XFILL_51_DFFSR_270 gnd vdd FILL
XFILL_75_DFFSR_32 gnd vdd FILL
XFILL_75_DFFSR_43 gnd vdd FILL
XFILL_15_3_1 gnd vdd FILL
XFILL_75_DFFSR_54 gnd vdd FILL
XFILL_75_DFFSR_65 gnd vdd FILL
XFILL_75_DFFSR_76 gnd vdd FILL
XFILL_75_DFFSR_87 gnd vdd FILL
XFILL_75_DFFSR_98 gnd vdd FILL
XFILL_3_INVX1_6 gnd vdd FILL
XFILL_10_NAND2X1_14 gnd vdd FILL
XFILL_10_NAND2X1_25 gnd vdd FILL
XFILL_44_DFFSR_20 gnd vdd FILL
XFILL_10_NAND2X1_36 gnd vdd FILL
XFILL_10_NAND2X1_47 gnd vdd FILL
XFILL_10_NAND2X1_58 gnd vdd FILL
XFILL_44_DFFSR_31 gnd vdd FILL
XFILL_10_NAND2X1_69 gnd vdd FILL
XFILL_15_NOR3X1_6 gnd vdd FILL
XFILL_44_DFFSR_42 gnd vdd FILL
XFILL_8_OAI22X1_19 gnd vdd FILL
XFILL_44_DFFSR_53 gnd vdd FILL
XFILL_44_DFFSR_64 gnd vdd FILL
XFILL_44_DFFSR_75 gnd vdd FILL
XFILL_82_DFFSR_180 gnd vdd FILL
XFILL_44_DFFSR_86 gnd vdd FILL
XFILL_82_DFFSR_191 gnd vdd FILL
XFILL_44_DFFSR_97 gnd vdd FILL
XFILL_33_DFFSR_204 gnd vdd FILL
XFILL_33_DFFSR_215 gnd vdd FILL
XFILL_84_DFFSR_30 gnd vdd FILL
XFILL_33_DFFSR_226 gnd vdd FILL
XFILL_33_DFFSR_237 gnd vdd FILL
XFILL_84_DFFSR_41 gnd vdd FILL
XFILL_2_DFFSR_250 gnd vdd FILL
XFILL_33_DFFSR_248 gnd vdd FILL
XFILL_84_DFFSR_52 gnd vdd FILL
XFILL_7_NAND3X1_40 gnd vdd FILL
XFILL_2_NAND3X1_110 gnd vdd FILL
XFILL_84_DFFSR_63 gnd vdd FILL
XFILL_2_NAND3X1_121 gnd vdd FILL
XFILL_2_DFFSR_261 gnd vdd FILL
XFILL_7_NAND3X1_51 gnd vdd FILL
XFILL_7_NAND3X1_62 gnd vdd FILL
XFILL_2_DFFSR_272 gnd vdd FILL
XFILL_2_NAND3X1_132 gnd vdd FILL
XFILL_84_DFFSR_74 gnd vdd FILL
XFILL_13_DFFSR_30 gnd vdd FILL
XFILL_33_DFFSR_259 gnd vdd FILL
XFILL_7_NAND3X1_73 gnd vdd FILL
XFILL_84_DFFSR_85 gnd vdd FILL
XFILL_86_DFFSR_190 gnd vdd FILL
XFILL_13_DFFSR_41 gnd vdd FILL
XFILL_60_DFFSR_104 gnd vdd FILL
XFILL_7_NAND3X1_84 gnd vdd FILL
XFILL_84_DFFSR_96 gnd vdd FILL
XFILL_37_DFFSR_203 gnd vdd FILL
XFILL_13_DFFSR_52 gnd vdd FILL
XFILL_13_DFFSR_63 gnd vdd FILL
XFILL_7_NAND3X1_95 gnd vdd FILL
XFILL_60_DFFSR_115 gnd vdd FILL
XFILL_13_DFFSR_74 gnd vdd FILL
XFILL_60_DFFSR_126 gnd vdd FILL
XFILL_37_DFFSR_214 gnd vdd FILL
XFILL_13_DFFSR_85 gnd vdd FILL
XFILL_37_DFFSR_225 gnd vdd FILL
XFILL_60_DFFSR_137 gnd vdd FILL
XFILL_37_DFFSR_236 gnd vdd FILL
XFILL_60_DFFSR_148 gnd vdd FILL
XFILL_13_DFFSR_96 gnd vdd FILL
XFILL_37_DFFSR_247 gnd vdd FILL
XFILL_6_DFFSR_260 gnd vdd FILL
XFILL_60_DFFSR_159 gnd vdd FILL
XFILL_6_DFFSR_271 gnd vdd FILL
XFILL_37_DFFSR_258 gnd vdd FILL
XFILL_53_DFFSR_40 gnd vdd FILL
XFILL_37_DFFSR_269 gnd vdd FILL
XFILL_3_MUX2X1_16 gnd vdd FILL
XFILL_24_NOR3X1_4 gnd vdd FILL
XFILL_3_MUX2X1_27 gnd vdd FILL
XFILL_53_DFFSR_51 gnd vdd FILL
XFILL_64_DFFSR_103 gnd vdd FILL
XFILL_64_DFFSR_114 gnd vdd FILL
XFILL_53_DFFSR_62 gnd vdd FILL
XFILL_3_MUX2X1_38 gnd vdd FILL
XFILL_19_CLKBUF1_17 gnd vdd FILL
XFILL_66_7_2 gnd vdd FILL
XFILL_19_CLKBUF1_28 gnd vdd FILL
XFILL_53_DFFSR_73 gnd vdd FILL
XFILL_3_MUX2X1_49 gnd vdd FILL
XFILL_64_DFFSR_125 gnd vdd FILL
XFILL_53_DFFSR_84 gnd vdd FILL
XFILL_19_CLKBUF1_39 gnd vdd FILL
XFILL_64_DFFSR_136 gnd vdd FILL
XFILL_53_DFFSR_95 gnd vdd FILL
XFILL_65_2_1 gnd vdd FILL
XFILL_14_AOI21X1_14 gnd vdd FILL
XFILL_64_DFFSR_147 gnd vdd FILL
XFILL_64_DFFSR_158 gnd vdd FILL
XFILL_14_AOI21X1_25 gnd vdd FILL
XFILL_14_AOI21X1_36 gnd vdd FILL
XFILL_64_DFFSR_169 gnd vdd FILL
XFILL_0_NAND2X1_20 gnd vdd FILL
XFILL_7_MUX2X1_15 gnd vdd FILL
XFILL_0_NAND2X1_31 gnd vdd FILL
XFILL_0_NAND2X1_42 gnd vdd FILL
XFILL_14_AOI21X1_47 gnd vdd FILL
XMUX2X1_40 INVX1_53/Y MUX2X1_7/B NAND2X1_5/Y gnd MUX2X1_40/Y vdd MUX2X1
XNOR2X1_101 DFFSR_159/Q NOR2X1_90/B gnd NOR2X1_101/Y vdd NOR2X1
XFILL_7_MUX2X1_26 gnd vdd FILL
XFILL_68_DFFSR_102 gnd vdd FILL
XMUX2X1_51 INVX1_64/Y BUFX4_65/Y NAND2X1_8/Y gnd MUX2X1_51/Y vdd MUX2X1
XFILL_0_NAND2X1_53 gnd vdd FILL
XFILL_7_MUX2X1_37 gnd vdd FILL
XNOR2X1_112 OAI21X1_46/B INVX1_163/Y gnd NAND2X1_6/B vdd NOR2X1
XFILL_14_AOI21X1_58 gnd vdd FILL
XFILL_14_AOI21X1_69 gnd vdd FILL
XNOR2X1_123 OR2X2_1/B INVX4_1/Y gnd AOI21X1_3/B vdd NOR2X1
XFILL_81_DFFSR_1 gnd vdd FILL
XFILL_68_DFFSR_113 gnd vdd FILL
XFILL_68_DFFSR_124 gnd vdd FILL
XFILL_7_MUX2X1_48 gnd vdd FILL
XMUX2X1_62 MUX2X1_66/A INVX1_75/Y NOR2X1_22/Y gnd MUX2X1_62/Y vdd MUX2X1
XFILL_0_NAND2X1_64 gnd vdd FILL
XMUX2X1_73 INVX1_86/Y BUFX4_64/Y OR2X2_1/Y gnd MUX2X1_73/Y vdd MUX2X1
XNOR2X1_134 DFFSR_142/Q AOI21X1_7/B gnd AOI21X1_7/C vdd NOR2X1
XFILL_68_DFFSR_135 gnd vdd FILL
XFILL_7_MUX2X1_59 gnd vdd FILL
XFILL_0_NAND2X1_75 gnd vdd FILL
XNOR2X1_145 DFFSR_104/Q AOI21X1_9/B gnd AOI21X1_9/C vdd NOR2X1
XMUX2X1_84 INVX1_97/Y BUFX4_64/Y MUX2X1_86/S gnd MUX2X1_84/Y vdd MUX2X1
XFILL_0_NAND2X1_86 gnd vdd FILL
XFILL_22_DFFSR_50 gnd vdd FILL
XFILL_68_DFFSR_146 gnd vdd FILL
XFILL_11_OAI21X1_3 gnd vdd FILL
XMUX2X1_95 MUX2X1_95/A BUFX4_96/Y MUX2X1_95/S gnd MUX2X1_95/Y vdd MUX2X1
XNOR2X1_156 NOR2X1_68/A NAND2X1_3/Y gnd NOR2X1_156/Y vdd NOR2X1
XFILL_68_DFFSR_157 gnd vdd FILL
XNOR2X1_167 NAND2X1_3/Y NOR2X1_10/B gnd NOR2X1_167/Y vdd NOR2X1
XFILL_22_DFFSR_61 gnd vdd FILL
XFILL_68_DFFSR_168 gnd vdd FILL
XNOR2X1_178 DFFSR_28/Q NOR2X1_181/B gnd NOR2X1_178/Y vdd NOR2X1
XFILL_22_DFFSR_72 gnd vdd FILL
XFILL_22_DFFSR_83 gnd vdd FILL
XFILL_68_DFFSR_179 gnd vdd FILL
XNOR2X1_189 DFFSR_21/Q NOR2X1_190/B gnd NOR2X1_189/Y vdd NOR2X1
XFILL_22_DFFSR_94 gnd vdd FILL
XFILL_7_NOR3X1_5 gnd vdd FILL
XFILL_15_OAI21X1_2 gnd vdd FILL
XFILL_62_DFFSR_60 gnd vdd FILL
XFILL_62_DFFSR_71 gnd vdd FILL
XFILL_62_DFFSR_82 gnd vdd FILL
XFILL_62_DFFSR_93 gnd vdd FILL
XFILL_3_INVX1_220 gnd vdd FILL
XFILL_26_CLKBUF1_30 gnd vdd FILL
XFILL_26_CLKBUF1_41 gnd vdd FILL
XFILL_5_DFFSR_40 gnd vdd FILL
XFILL_46_DFFSR_4 gnd vdd FILL
XFILL_5_DFFSR_51 gnd vdd FILL
XFILL_9_CLKBUF1_12 gnd vdd FILL
XFILL_5_DFFSR_62 gnd vdd FILL
XMUX2X1_107 BUFX4_78/Y INVX1_1/Y MUX2X1_1/S gnd DFFSR_185/D vdd MUX2X1
XMUX2X1_118 MUX2X1_2/A INVX1_112/Y MUX2X1_1/S gnd DFFSR_186/D vdd MUX2X1
XFILL_5_DFFSR_73 gnd vdd FILL
XFILL_5_DFFSR_84 gnd vdd FILL
XMUX2X1_129 BUFX4_87/Y NOR3X1_49/A AOI21X1_1/B gnd DFFSR_178/D vdd MUX2X1
XFILL_9_CLKBUF1_23 gnd vdd FILL
XFILL_23_MUX2X1_13 gnd vdd FILL
XFILL_5_DFFSR_95 gnd vdd FILL
XFILL_9_CLKBUF1_34 gnd vdd FILL
XFILL_31_DFFSR_70 gnd vdd FILL
XFILL_23_MUX2X1_24 gnd vdd FILL
XFILL_23_MUX2X1_35 gnd vdd FILL
XFILL_31_DFFSR_81 gnd vdd FILL
XFILL_17_MUX2X1_108 gnd vdd FILL
XFILL_17_MUX2X1_119 gnd vdd FILL
XFILL_31_DFFSR_92 gnd vdd FILL
XFILL_4_AOI21X1_20 gnd vdd FILL
XFILL_23_MUX2X1_46 gnd vdd FILL
XFILL_4_AOI21X1_31 gnd vdd FILL
XFILL_23_MUX2X1_57 gnd vdd FILL
XFILL_4_AOI21X1_42 gnd vdd FILL
XFILL_23_MUX2X1_68 gnd vdd FILL
XFILL_23_MUX2X1_79 gnd vdd FILL
XFILL_4_AOI21X1_53 gnd vdd FILL
XFILL_14_OAI22X1_11 gnd vdd FILL
XFILL_14_OAI22X1_22 gnd vdd FILL
XFILL_4_AOI21X1_64 gnd vdd FILL
XFILL_9_BUFX2_9 gnd vdd FILL
XFILL_53_DFFSR_190 gnd vdd FILL
XFILL_4_AOI21X1_75 gnd vdd FILL
XFILL_14_OAI22X1_33 gnd vdd FILL
XINVX1_14 INVX1_14/A gnd INVX1_14/Y vdd INVX1
XFILL_71_DFFSR_80 gnd vdd FILL
XFILL_14_OAI22X1_44 gnd vdd FILL
XINVX1_25 INVX1_25/A gnd NOR3X1_4/A vdd INVX1
XINVX1_36 DFFSR_4/Q gnd INVX1_36/Y vdd INVX1
XFILL_71_DFFSR_91 gnd vdd FILL
XINVX1_47 INVX1_47/A gnd INVX1_47/Y vdd INVX1
XFILL_7_NOR2X1_130 gnd vdd FILL
XFILL_7_NOR2X1_141 gnd vdd FILL
XINVX1_58 INVX1_58/A gnd INVX1_58/Y vdd INVX1
XINVX1_69 INVX1_69/A gnd INVX1_69/Y vdd INVX1
XFILL_57_7_2 gnd vdd FILL
XFILL_7_NOR2X1_152 gnd vdd FILL
XFILL_7_NOR2X1_163 gnd vdd FILL
XFILL_7_NOR2X1_174 gnd vdd FILL
XFILL_56_2_1 gnd vdd FILL
XFILL_31_DFFSR_103 gnd vdd FILL
XFILL_7_NOR2X1_185 gnd vdd FILL
XFILL_31_DFFSR_114 gnd vdd FILL
XFILL_7_NOR2X1_196 gnd vdd FILL
XFILL_68_DFFSR_8 gnd vdd FILL
XFILL_31_DFFSR_125 gnd vdd FILL
XFILL_31_DFFSR_136 gnd vdd FILL
XFILL_0_DFFSR_160 gnd vdd FILL
XFILL_11_NOR2X1_202 gnd vdd FILL
XFILL_31_DFFSR_147 gnd vdd FILL
XFILL_31_DFFSR_158 gnd vdd FILL
XFILL_0_DFFSR_171 gnd vdd FILL
XFILL_40_DFFSR_90 gnd vdd FILL
XFILL_31_DFFSR_169 gnd vdd FILL
XFILL_0_DFFSR_182 gnd vdd FILL
XFILL_0_DFFSR_193 gnd vdd FILL
XFILL_35_DFFSR_102 gnd vdd FILL
XFILL_35_DFFSR_113 gnd vdd FILL
XFILL_35_DFFSR_124 gnd vdd FILL
XFILL_35_DFFSR_135 gnd vdd FILL
XFILL_35_DFFSR_146 gnd vdd FILL
XFILL_35_DFFSR_157 gnd vdd FILL
XFILL_4_DFFSR_170 gnd vdd FILL
XFILL_35_DFFSR_168 gnd vdd FILL
XFILL_4_DFFSR_181 gnd vdd FILL
XFILL_35_DFFSR_179 gnd vdd FILL
XFILL_40_6_2 gnd vdd FILL
XFILL_4_DFFSR_192 gnd vdd FILL
XFILL_7_MUX2X1_103 gnd vdd FILL
XFILL_39_DFFSR_101 gnd vdd FILL
XFILL_7_MUX2X1_114 gnd vdd FILL
XFILL_39_DFFSR_112 gnd vdd FILL
XFILL_7_MUX2X1_125 gnd vdd FILL
XFILL_39_DFFSR_123 gnd vdd FILL
XFILL_39_DFFSR_134 gnd vdd FILL
XFILL_7_MUX2X1_136 gnd vdd FILL
XFILL_8_BUFX4_3 gnd vdd FILL
XFILL_39_DFFSR_145 gnd vdd FILL
XFILL_7_MUX2X1_147 gnd vdd FILL
XFILL_7_MUX2X1_158 gnd vdd FILL
XFILL_39_DFFSR_156 gnd vdd FILL
XFILL_8_DFFSR_180 gnd vdd FILL
XFILL_39_DFFSR_167 gnd vdd FILL
XFILL_7_MUX2X1_169 gnd vdd FILL
XFILL_39_DFFSR_178 gnd vdd FILL
XFILL_8_DFFSR_191 gnd vdd FILL
XFILL_31_NOR3X1_14 gnd vdd FILL
XFILL_4_OAI22X1_50 gnd vdd FILL
XFILL_39_DFFSR_189 gnd vdd FILL
XFILL_31_NOR3X1_25 gnd vdd FILL
XFILL_31_NOR3X1_36 gnd vdd FILL
XFILL_8_OAI21X1_30 gnd vdd FILL
XFILL_31_NOR3X1_47 gnd vdd FILL
XFILL_81_DFFSR_203 gnd vdd FILL
XFILL_8_OAI21X1_41 gnd vdd FILL
XFILL_81_DFFSR_214 gnd vdd FILL
XFILL_81_DFFSR_225 gnd vdd FILL
XFILL_81_DFFSR_236 gnd vdd FILL
XFILL_81_DFFSR_247 gnd vdd FILL
XFILL_81_DFFSR_258 gnd vdd FILL
XFILL_81_DFFSR_269 gnd vdd FILL
XFILL_85_DFFSR_202 gnd vdd FILL
XFILL_85_DFFSR_213 gnd vdd FILL
XFILL_85_DFFSR_224 gnd vdd FILL
XFILL_85_DFFSR_235 gnd vdd FILL
XFILL_12_AOI21X1_9 gnd vdd FILL
XFILL_85_DFFSR_246 gnd vdd FILL
XFILL_7_INVX1_7 gnd vdd FILL
XFILL_85_DFFSR_257 gnd vdd FILL
XFILL_85_DFFSR_268 gnd vdd FILL
XFILL_20_DFFSR_190 gnd vdd FILL
XFILL_1_INVX1_130 gnd vdd FILL
XFILL_48_7_2 gnd vdd FILL
XFILL_1_INVX1_141 gnd vdd FILL
XFILL_1_INVX1_152 gnd vdd FILL
XFILL_1_INVX1_163 gnd vdd FILL
XFILL_47_2_1 gnd vdd FILL
XFILL_1_INVX1_174 gnd vdd FILL
XFILL_1_INVX1_185 gnd vdd FILL
XFILL_8_NAND3X1_104 gnd vdd FILL
XFILL_8_NAND3X1_115 gnd vdd FILL
XFILL_8_NAND3X1_126 gnd vdd FILL
XFILL_1_INVX1_196 gnd vdd FILL
XFILL_5_INVX1_140 gnd vdd FILL
XFILL_5_INVX1_151 gnd vdd FILL
XFILL_5_INVX1_162 gnd vdd FILL
XFILL_5_INVX1_173 gnd vdd FILL
XFILL_5_INVX1_184 gnd vdd FILL
XFILL_5_INVX1_195 gnd vdd FILL
XFILL_31_6_2 gnd vdd FILL
XFILL_30_1_1 gnd vdd FILL
XFILL_3_OAI22X1_2 gnd vdd FILL
XFILL_3_NAND2X1_19 gnd vdd FILL
XFILL_28_DFFSR_1 gnd vdd FILL
XFILL_85_DFFSR_2 gnd vdd FILL
XFILL_7_OAI22X1_1 gnd vdd FILL
XFILL_3_NAND3X1_100 gnd vdd FILL
XFILL_3_NAND3X1_111 gnd vdd FILL
XFILL_13_MUX2X1_150 gnd vdd FILL
XFILL_3_NAND3X1_122 gnd vdd FILL
XFILL_13_MUX2X1_161 gnd vdd FILL
XFILL_13_MUX2X1_172 gnd vdd FILL
XFILL_13_MUX2X1_183 gnd vdd FILL
XFILL_52_DFFSR_202 gnd vdd FILL
XFILL_13_MUX2X1_194 gnd vdd FILL
XFILL_52_DFFSR_213 gnd vdd FILL
XFILL_52_DFFSR_224 gnd vdd FILL
XFILL_52_DFFSR_235 gnd vdd FILL
XFILL_52_DFFSR_246 gnd vdd FILL
XFILL_85_DFFSR_19 gnd vdd FILL
XFILL_39_7_2 gnd vdd FILL
XFILL_52_DFFSR_257 gnd vdd FILL
XFILL_52_DFFSR_268 gnd vdd FILL
XFILL_12_DFFSR_7 gnd vdd FILL
XFILL_56_DFFSR_201 gnd vdd FILL
XFILL_38_2_1 gnd vdd FILL
XFILL_14_DFFSR_19 gnd vdd FILL
XFILL_29_CLKBUF1_18 gnd vdd FILL
XFILL_29_CLKBUF1_29 gnd vdd FILL
XFILL_56_DFFSR_212 gnd vdd FILL
XFILL_56_DFFSR_223 gnd vdd FILL
XFILL_56_DFFSR_234 gnd vdd FILL
XFILL_56_DFFSR_245 gnd vdd FILL
XFILL_56_DFFSR_256 gnd vdd FILL
XFILL_56_DFFSR_267 gnd vdd FILL
XFILL_11_CLKBUF1_8 gnd vdd FILL
XFILL_83_DFFSR_101 gnd vdd FILL
XFILL_54_DFFSR_18 gnd vdd FILL
XFILL_83_DFFSR_112 gnd vdd FILL
XFILL_54_DFFSR_29 gnd vdd FILL
XFILL_83_DFFSR_123 gnd vdd FILL
XFILL_83_DFFSR_134 gnd vdd FILL
XFILL_7_AOI21X1_19 gnd vdd FILL
XFILL_83_DFFSR_145 gnd vdd FILL
XFILL_83_DFFSR_156 gnd vdd FILL
XFILL_83_DFFSR_167 gnd vdd FILL
XFILL_22_6_2 gnd vdd FILL
XFILL_15_CLKBUF1_7 gnd vdd FILL
XFILL_83_DFFSR_178 gnd vdd FILL
XFILL_83_DFFSR_189 gnd vdd FILL
XFILL_87_DFFSR_100 gnd vdd FILL
XFILL_21_1_1 gnd vdd FILL
XFILL_3_DFFSR_204 gnd vdd FILL
XFILL_0_NAND3X1_4 gnd vdd FILL
XFILL_3_DFFSR_215 gnd vdd FILL
XFILL_87_DFFSR_111 gnd vdd FILL
XFILL_3_DFFSR_226 gnd vdd FILL
XFILL_87_DFFSR_122 gnd vdd FILL
XFILL_87_DFFSR_133 gnd vdd FILL
XFILL_3_DFFSR_237 gnd vdd FILL
XFILL_87_DFFSR_144 gnd vdd FILL
XFILL_3_DFFSR_248 gnd vdd FILL
XFILL_87_DFFSR_155 gnd vdd FILL
XFILL_11_BUFX4_102 gnd vdd FILL
XFILL_23_DFFSR_17 gnd vdd FILL
XFILL_3_DFFSR_259 gnd vdd FILL
XFILL_23_DFFSR_28 gnd vdd FILL
XFILL_87_DFFSR_166 gnd vdd FILL
XFILL_87_DFFSR_177 gnd vdd FILL
XFILL_14_BUFX4_60 gnd vdd FILL
XFILL_23_DFFSR_39 gnd vdd FILL
XFILL_19_CLKBUF1_6 gnd vdd FILL
XFILL_14_BUFX4_71 gnd vdd FILL
XFILL_87_DFFSR_188 gnd vdd FILL
XFILL_7_DFFSR_203 gnd vdd FILL
XFILL_4_NAND3X1_3 gnd vdd FILL
XFILL_87_DFFSR_199 gnd vdd FILL
XFILL_7_DFFSR_214 gnd vdd FILL
XFILL_14_BUFX4_82 gnd vdd FILL
XFILL_14_BUFX4_93 gnd vdd FILL
XFILL_7_DFFSR_225 gnd vdd FILL
XFILL_7_DFFSR_236 gnd vdd FILL
XDFFSR_250 INVX1_47/A CLKBUF1_5/Y BUFX4_50/Y vdd MUX2X1_33/Y gnd vdd DFFSR
XFILL_7_DFFSR_247 gnd vdd FILL
XDFFSR_261 NOR2X1_16/A DFFSR_5/CLK DFFSR_5/R vdd DFFSR_261/D gnd vdd DFFSR
XDFFSR_272 NOR2X1_4/A DFFSR_8/CLK DFFSR_8/R vdd DFFSR_272/D gnd vdd DFFSR
XFILL_7_DFFSR_258 gnd vdd FILL
XFILL_15_BUFX4_101 gnd vdd FILL
XFILL_63_DFFSR_16 gnd vdd FILL
XFILL_7_DFFSR_269 gnd vdd FILL
XFILL_63_DFFSR_27 gnd vdd FILL
XFILL_63_DFFSR_38 gnd vdd FILL
XFILL_63_DFFSR_49 gnd vdd FILL
XFILL_8_NAND3X1_2 gnd vdd FILL
XFILL_6_DFFSR_18 gnd vdd FILL
XFILL_6_DFFSR_29 gnd vdd FILL
XFILL_32_DFFSR_15 gnd vdd FILL
XFILL_32_DFFSR_26 gnd vdd FILL
XFILL_32_DFFSR_37 gnd vdd FILL
XFILL_5_7_2 gnd vdd FILL
XFILL_32_DFFSR_48 gnd vdd FILL
XFILL_0_AOI22X1_9 gnd vdd FILL
XFILL_32_DFFSR_59 gnd vdd FILL
XFILL_7_OAI22X1_16 gnd vdd FILL
XFILL_29_2_1 gnd vdd FILL
XFILL_4_2_1 gnd vdd FILL
XFILL_7_OAI22X1_27 gnd vdd FILL
XFILL_7_OAI22X1_38 gnd vdd FILL
XFILL_7_OAI22X1_49 gnd vdd FILL
XFILL_72_DFFSR_14 gnd vdd FILL
XFILL_23_DFFSR_201 gnd vdd FILL
XFILL_0_INVX1_208 gnd vdd FILL
XFILL_72_DFFSR_25 gnd vdd FILL
XFILL_0_INVX1_219 gnd vdd FILL
XFILL_72_DFFSR_36 gnd vdd FILL
XFILL_23_DFFSR_212 gnd vdd FILL
XFILL_23_DFFSR_223 gnd vdd FILL
XFILL_72_DFFSR_47 gnd vdd FILL
XFILL_23_DFFSR_234 gnd vdd FILL
XFILL_72_DFFSR_58 gnd vdd FILL
XFILL_15_MUX2X1_4 gnd vdd FILL
XFILL_4_AOI22X1_8 gnd vdd FILL
XFILL_72_DFFSR_69 gnd vdd FILL
XFILL_23_DFFSR_245 gnd vdd FILL
XFILL_23_DFFSR_256 gnd vdd FILL
XFILL_23_DFFSR_267 gnd vdd FILL
XFILL_6_NAND3X1_70 gnd vdd FILL
XFILL_6_NAND3X1_81 gnd vdd FILL
XFILL_4_INVX1_207 gnd vdd FILL
XFILL_50_DFFSR_101 gnd vdd FILL
XFILL_27_DFFSR_200 gnd vdd FILL
XFILL_27_DFFSR_211 gnd vdd FILL
XFILL_6_NAND3X1_92 gnd vdd FILL
XFILL_50_DFFSR_112 gnd vdd FILL
XFILL_4_INVX1_218 gnd vdd FILL
XFILL_50_DFFSR_123 gnd vdd FILL
XFILL_50_DFFSR_134 gnd vdd FILL
XFILL_27_DFFSR_222 gnd vdd FILL
XFILL_13_6_2 gnd vdd FILL
XFILL_8_AOI22X1_7 gnd vdd FILL
XFILL_41_DFFSR_13 gnd vdd FILL
XFILL_27_DFFSR_233 gnd vdd FILL
XFILL_6_BUFX4_70 gnd vdd FILL
XFILL_41_DFFSR_24 gnd vdd FILL
XFILL_50_DFFSR_145 gnd vdd FILL
XFILL_27_DFFSR_244 gnd vdd FILL
XFILL_50_DFFSR_156 gnd vdd FILL
XFILL_6_BUFX4_81 gnd vdd FILL
XFILL_27_DFFSR_255 gnd vdd FILL
XFILL_12_1_1 gnd vdd FILL
XFILL_41_DFFSR_35 gnd vdd FILL
XFILL_6_BUFX4_92 gnd vdd FILL
XFILL_50_DFFSR_167 gnd vdd FILL
XFILL_50_DFFSR_178 gnd vdd FILL
XFILL_41_DFFSR_46 gnd vdd FILL
XFILL_27_DFFSR_266 gnd vdd FILL
XFILL_41_DFFSR_57 gnd vdd FILL
XFILL_0_OAI21X1_18 gnd vdd FILL
XFILL_0_OAI21X1_29 gnd vdd FILL
XFILL_41_DFFSR_68 gnd vdd FILL
XFILL_54_DFFSR_100 gnd vdd FILL
XFILL_50_DFFSR_189 gnd vdd FILL
XFILL_54_DFFSR_111 gnd vdd FILL
XFILL_41_DFFSR_79 gnd vdd FILL
XFILL_18_CLKBUF1_14 gnd vdd FILL
XFILL_18_CLKBUF1_25 gnd vdd FILL
XFILL_54_DFFSR_122 gnd vdd FILL
XFILL_18_CLKBUF1_36 gnd vdd FILL
XFILL_54_DFFSR_133 gnd vdd FILL
XFILL_81_DFFSR_12 gnd vdd FILL
XFILL_13_AOI21X1_11 gnd vdd FILL
XFILL_54_DFFSR_144 gnd vdd FILL
XFILL_81_DFFSR_23 gnd vdd FILL
XFILL_54_DFFSR_155 gnd vdd FILL
XFILL_13_AOI21X1_22 gnd vdd FILL
XFILL_81_DFFSR_34 gnd vdd FILL
XFILL_13_AOI21X1_33 gnd vdd FILL
XFILL_54_DFFSR_166 gnd vdd FILL
XFILL_54_DFFSR_177 gnd vdd FILL
XFILL_81_DFFSR_45 gnd vdd FILL
XFILL_13_AOI21X1_44 gnd vdd FILL
XFILL_81_DFFSR_56 gnd vdd FILL
XFILL_10_DFFSR_12 gnd vdd FILL
XFILL_54_DFFSR_188 gnd vdd FILL
XFILL_81_DFFSR_67 gnd vdd FILL
XFILL_10_DFFSR_23 gnd vdd FILL
XFILL_13_AOI21X1_55 gnd vdd FILL
XFILL_13_AOI21X1_66 gnd vdd FILL
XFILL_81_DFFSR_78 gnd vdd FILL
XFILL_10_DFFSR_34 gnd vdd FILL
XFILL_58_DFFSR_110 gnd vdd FILL
XFILL_54_DFFSR_199 gnd vdd FILL
XFILL_81_DFFSR_89 gnd vdd FILL
XFILL_13_AOI21X1_77 gnd vdd FILL
XFILL_58_DFFSR_121 gnd vdd FILL
XFILL_58_DFFSR_132 gnd vdd FILL
XFILL_10_DFFSR_45 gnd vdd FILL
XFILL_10_DFFSR_56 gnd vdd FILL
XFILL_58_DFFSR_143 gnd vdd FILL
XFILL_10_DFFSR_67 gnd vdd FILL
XFILL_8_NOR2X1_5 gnd vdd FILL
XFILL_58_DFFSR_154 gnd vdd FILL
XFILL_10_DFFSR_78 gnd vdd FILL
XFILL_10_DFFSR_89 gnd vdd FILL
XFILL_58_DFFSR_165 gnd vdd FILL
XFILL_58_DFFSR_176 gnd vdd FILL
XFILL_50_DFFSR_11 gnd vdd FILL
XFILL_1_DFFSR_103 gnd vdd FILL
XFILL_58_DFFSR_187 gnd vdd FILL
XFILL_58_DFFSR_198 gnd vdd FILL
XFILL_50_DFFSR_22 gnd vdd FILL
XFILL_1_DFFSR_114 gnd vdd FILL
XFILL_50_DFFSR_33 gnd vdd FILL
XFILL_1_DFFSR_125 gnd vdd FILL
XFILL_1_DFFSR_136 gnd vdd FILL
XFILL_21_NOR3X1_8 gnd vdd FILL
XFILL_50_DFFSR_44 gnd vdd FILL
XFILL_8_5 gnd vdd FILL
XFILL_50_DFFSR_55 gnd vdd FILL
XFILL_1_DFFSR_147 gnd vdd FILL
XFILL_1_DFFSR_158 gnd vdd FILL
XFILL_50_DFFSR_66 gnd vdd FILL
XFILL_50_DFFSR_77 gnd vdd FILL
XFILL_1_DFFSR_169 gnd vdd FILL
XFILL_50_DFFSR_88 gnd vdd FILL
XFILL_50_DFFSR_99 gnd vdd FILL
XFILL_5_DFFSR_102 gnd vdd FILL
XFILL_7_MUX2X1_3 gnd vdd FILL
XFILL_5_DFFSR_113 gnd vdd FILL
XFILL_5_DFFSR_124 gnd vdd FILL
XFILL_5_DFFSR_135 gnd vdd FILL
XFILL_5_DFFSR_146 gnd vdd FILL
XFILL_5_DFFSR_157 gnd vdd FILL
XFILL_51_DFFSR_5 gnd vdd FILL
XFILL_5_DFFSR_168 gnd vdd FILL
XFILL_5_DFFSR_179 gnd vdd FILL
XFILL_9_NAND3X1_105 gnd vdd FILL
XFILL_63_5_2 gnd vdd FILL
XFILL_8_CLKBUF1_20 gnd vdd FILL
XFILL_9_DFFSR_101 gnd vdd FILL
XFILL_9_NAND3X1_116 gnd vdd FILL
XFILL_13_MUX2X1_10 gnd vdd FILL
XFILL_9_NAND3X1_127 gnd vdd FILL
XFILL_9_DFFSR_112 gnd vdd FILL
XFILL_13_MUX2X1_21 gnd vdd FILL
XFILL_8_CLKBUF1_31 gnd vdd FILL
XFILL_9_DFFSR_123 gnd vdd FILL
XFILL_9_DFFSR_134 gnd vdd FILL
XFILL_62_0_1 gnd vdd FILL
XFILL_13_MUX2X1_32 gnd vdd FILL
XFILL_8_CLKBUF1_42 gnd vdd FILL
XFILL_9_DFFSR_145 gnd vdd FILL
XFILL_16_MUX2X1_105 gnd vdd FILL
XFILL_13_MUX2X1_43 gnd vdd FILL
XFILL_4_NOR3X1_9 gnd vdd FILL
XFILL_16_MUX2X1_116 gnd vdd FILL
XFILL_9_DFFSR_156 gnd vdd FILL
XFILL_13_MUX2X1_54 gnd vdd FILL
XFILL_16_MUX2X1_127 gnd vdd FILL
XFILL_9_DFFSR_167 gnd vdd FILL
XFILL_16_MUX2X1_138 gnd vdd FILL
XFILL_13_MUX2X1_65 gnd vdd FILL
XFILL_9_DFFSR_178 gnd vdd FILL
XFILL_1_NOR3X1_14 gnd vdd FILL
XFILL_13_MUX2X1_76 gnd vdd FILL
XFILL_3_AOI21X1_50 gnd vdd FILL
XFILL_30_NOR3X1_6 gnd vdd FILL
XFILL_13_MUX2X1_87 gnd vdd FILL
XFILL_16_MUX2X1_149 gnd vdd FILL
XFILL_9_DFFSR_189 gnd vdd FILL
XFILL_3_AOI21X1_61 gnd vdd FILL
XOAI21X1_20 INVX1_168/Y OAI21X1_2/B OAI21X1_20/C gnd NOR2X1_92/B vdd OAI21X1
XFILL_1_NOR3X1_25 gnd vdd FILL
XFILL_3_AOI21X1_72 gnd vdd FILL
XFILL_1_NOR3X1_36 gnd vdd FILL
XOAI21X1_31 INVX1_195/Y OAI21X1_6/B OAI21X1_31/C gnd OAI21X1_31/Y vdd OAI21X1
XFILL_13_OAI22X1_30 gnd vdd FILL
XFILL_13_MUX2X1_98 gnd vdd FILL
XFILL_13_OAI22X1_41 gnd vdd FILL
XFILL_1_NOR3X1_47 gnd vdd FILL
XFILL_17_MUX2X1_20 gnd vdd FILL
XFILL_17_MUX2X1_31 gnd vdd FILL
XOAI21X1_42 OAI21X1_45/A OAI21X1_45/B INVX2_5/Y gnd OAI21X1_42/Y vdd OAI21X1
XFILL_17_MUX2X1_42 gnd vdd FILL
XFILL_17_MUX2X1_53 gnd vdd FILL
XFILL_17_MUX2X1_64 gnd vdd FILL
XFILL_2_DFFSR_11 gnd vdd FILL
XFILL_5_NOR3X1_13 gnd vdd FILL
XFILL_17_MUX2X1_75 gnd vdd FILL
XFILL_2_DFFSR_22 gnd vdd FILL
XFILL_17_MUX2X1_86 gnd vdd FILL
XFILL_2_DFFSR_33 gnd vdd FILL
XFILL_6_NOR2X1_160 gnd vdd FILL
XFILL_17_MUX2X1_97 gnd vdd FILL
XFILL_5_NOR3X1_24 gnd vdd FILL
XFILL_2_DFFSR_44 gnd vdd FILL
XFILL_2_DFFSR_55 gnd vdd FILL
XFILL_5_NOR3X1_35 gnd vdd FILL
XFILL_16_DFFSR_8 gnd vdd FILL
XFILL_6_NOR2X1_171 gnd vdd FILL
XFILL_5_NOR3X1_46 gnd vdd FILL
XFILL_21_DFFSR_100 gnd vdd FILL
XFILL_6_NOR2X1_182 gnd vdd FILL
XFILL_73_DFFSR_9 gnd vdd FILL
XFILL_6_NOR2X1_193 gnd vdd FILL
XFILL_2_DFFSR_66 gnd vdd FILL
XFILL_21_DFFSR_111 gnd vdd FILL
XFILL_2_DFFSR_77 gnd vdd FILL
XFILL_21_DFFSR_122 gnd vdd FILL
XFILL_21_DFFSR_133 gnd vdd FILL
XFILL_2_DFFSR_88 gnd vdd FILL
XFILL_2_DFFSR_99 gnd vdd FILL
XFILL_21_DFFSR_144 gnd vdd FILL
XFILL_21_DFFSR_155 gnd vdd FILL
XFILL_9_NOR3X1_12 gnd vdd FILL
XFILL_9_NOR3X1_23 gnd vdd FILL
XFILL_21_DFFSR_166 gnd vdd FILL
XFILL_21_DFFSR_177 gnd vdd FILL
XFILL_9_NOR3X1_34 gnd vdd FILL
XFILL_2_INVX1_106 gnd vdd FILL
XFILL_21_DFFSR_188 gnd vdd FILL
XFILL_2_INVX1_117 gnd vdd FILL
XFILL_9_NOR3X1_45 gnd vdd FILL
XFILL_2_INVX1_128 gnd vdd FILL
XFILL_25_DFFSR_110 gnd vdd FILL
XFILL_21_DFFSR_199 gnd vdd FILL
XFILL_25_DFFSR_121 gnd vdd FILL
XFILL_25_DFFSR_132 gnd vdd FILL
XFILL_2_INVX1_139 gnd vdd FILL
XFILL_25_DFFSR_143 gnd vdd FILL
XFILL_25_DFFSR_154 gnd vdd FILL
XFILL_23_MUX2X1_140 gnd vdd FILL
XFILL_4_NAND3X1_101 gnd vdd FILL
XFILL_25_DFFSR_165 gnd vdd FILL
XFILL_4_NAND3X1_112 gnd vdd FILL
XFILL_4_NAND3X1_123 gnd vdd FILL
XFILL_25_DFFSR_176 gnd vdd FILL
XFILL_23_MUX2X1_151 gnd vdd FILL
XFILL_6_MUX2X1_100 gnd vdd FILL
XFILL_6_INVX1_105 gnd vdd FILL
XFILL_23_MUX2X1_162 gnd vdd FILL
XFILL_25_DFFSR_187 gnd vdd FILL
XFILL_6_MUX2X1_111 gnd vdd FILL
XFILL_23_MUX2X1_173 gnd vdd FILL
XFILL_6_INVX1_116 gnd vdd FILL
XFILL_6_INVX1_127 gnd vdd FILL
XFILL_25_DFFSR_198 gnd vdd FILL
XFILL_23_MUX2X1_184 gnd vdd FILL
XFILL_6_MUX2X1_122 gnd vdd FILL
XFILL_29_DFFSR_120 gnd vdd FILL
XFILL_6_INVX1_138 gnd vdd FILL
XFILL_29_DFFSR_131 gnd vdd FILL
XFILL_6_MUX2X1_133 gnd vdd FILL
XFILL_6_MUX2X1_144 gnd vdd FILL
XFILL_29_DFFSR_142 gnd vdd FILL
XFILL_6_INVX1_149 gnd vdd FILL
XFILL_6_MUX2X1_155 gnd vdd FILL
XFILL_29_DFFSR_153 gnd vdd FILL
XFILL_6_MUX2X1_166 gnd vdd FILL
XFILL_29_DFFSR_164 gnd vdd FILL
XFILL_21_NOR3X1_11 gnd vdd FILL
XFILL_29_DFFSR_175 gnd vdd FILL
XFILL_6_MUX2X1_177 gnd vdd FILL
XFILL_29_DFFSR_186 gnd vdd FILL
XFILL_6_MUX2X1_188 gnd vdd FILL
XFILL_29_DFFSR_197 gnd vdd FILL
XFILL_21_NOR3X1_22 gnd vdd FILL
XFILL_21_NOR3X1_33 gnd vdd FILL
XFILL_71_DFFSR_200 gnd vdd FILL
XFILL_21_NOR3X1_44 gnd vdd FILL
XFILL_71_DFFSR_211 gnd vdd FILL
XFILL_54_5_2 gnd vdd FILL
XFILL_71_DFFSR_222 gnd vdd FILL
XFILL_71_DFFSR_233 gnd vdd FILL
XFILL_53_0_1 gnd vdd FILL
XFILL_71_DFFSR_244 gnd vdd FILL
XFILL_25_NOR3X1_10 gnd vdd FILL
XFILL_71_DFFSR_255 gnd vdd FILL
XFILL_25_NOR3X1_21 gnd vdd FILL
XFILL_71_DFFSR_266 gnd vdd FILL
XFILL_25_NOR3X1_32 gnd vdd FILL
XFILL_25_NOR3X1_43 gnd vdd FILL
XFILL_75_DFFSR_210 gnd vdd FILL
XFILL_75_DFFSR_221 gnd vdd FILL
XFILL_75_DFFSR_232 gnd vdd FILL
XFILL_75_DFFSR_243 gnd vdd FILL
XFILL_10_BUFX4_8 gnd vdd FILL
XFILL_75_DFFSR_254 gnd vdd FILL
XFILL_75_DFFSR_265 gnd vdd FILL
XFILL_29_NOR3X1_20 gnd vdd FILL
XFILL_29_NOR3X1_31 gnd vdd FILL
XFILL_30_CLKBUF1_6 gnd vdd FILL
XFILL_29_NOR3X1_42 gnd vdd FILL
XFILL_79_DFFSR_220 gnd vdd FILL
XFILL_79_DFFSR_231 gnd vdd FILL
XFILL_79_DFFSR_242 gnd vdd FILL
XFILL_79_DFFSR_253 gnd vdd FILL
XFILL_79_DFFSR_264 gnd vdd FILL
XFILL_79_DFFSR_275 gnd vdd FILL
XFILL_34_CLKBUF1_5 gnd vdd FILL
XFILL_9_NAND3X1_14 gnd vdd FILL
XFILL_9_NAND3X1_25 gnd vdd FILL
XFILL_9_NAND3X1_36 gnd vdd FILL
XFILL_9_NAND3X1_47 gnd vdd FILL
XFILL_9_NAND3X1_58 gnd vdd FILL
XFILL_9_NAND3X1_69 gnd vdd FILL
XFILL_15_BUFX4_16 gnd vdd FILL
XFILL_15_BUFX4_27 gnd vdd FILL
XFILL_0_NOR3X1_2 gnd vdd FILL
XFILL_15_BUFX4_38 gnd vdd FILL
XFILL_15_BUFX4_49 gnd vdd FILL
XFILL_2_NAND2X1_16 gnd vdd FILL
XFILL_33_DFFSR_2 gnd vdd FILL
XFILL_2_NAND2X1_27 gnd vdd FILL
XFILL_45_5_2 gnd vdd FILL
XFILL_2_NAND2X1_38 gnd vdd FILL
XFILL_2_NAND2X1_49 gnd vdd FILL
XFILL_44_0_1 gnd vdd FILL
XFILL_0_OAI21X1_1 gnd vdd FILL
XFILL_12_MUX2X1_180 gnd vdd FILL
XFILL_12_MUX2X1_191 gnd vdd FILL
XFILL_42_DFFSR_210 gnd vdd FILL
XFILL_42_DFFSR_221 gnd vdd FILL
XFILL_42_DFFSR_232 gnd vdd FILL
XFILL_42_DFFSR_243 gnd vdd FILL
XFILL_42_DFFSR_254 gnd vdd FILL
XFILL_1_NOR2X1_80 gnd vdd FILL
XFILL_42_DFFSR_265 gnd vdd FILL
XFILL_1_NOR2X1_91 gnd vdd FILL
XFILL_28_CLKBUF1_15 gnd vdd FILL
XFILL_28_CLKBUF1_26 gnd vdd FILL
XFILL_55_DFFSR_6 gnd vdd FILL
XFILL_46_DFFSR_220 gnd vdd FILL
XFILL_28_CLKBUF1_37 gnd vdd FILL
XFILL_7_BUFX4_15 gnd vdd FILL
XFILL_46_DFFSR_231 gnd vdd FILL
XFILL_46_DFFSR_242 gnd vdd FILL
XFILL_7_BUFX4_26 gnd vdd FILL
XFILL_46_DFFSR_253 gnd vdd FILL
XFILL_7_BUFX4_37 gnd vdd FILL
XFILL_46_DFFSR_264 gnd vdd FILL
XFILL_7_BUFX4_48 gnd vdd FILL
XFILL_46_DFFSR_275 gnd vdd FILL
XFILL_5_NOR2X1_90 gnd vdd FILL
XFILL_7_BUFX4_59 gnd vdd FILL
XFILL_73_DFFSR_120 gnd vdd FILL
XFILL_73_DFFSR_131 gnd vdd FILL
XFILL_6_AOI21X1_16 gnd vdd FILL
XFILL_73_DFFSR_142 gnd vdd FILL
XFILL_6_AOI21X1_27 gnd vdd FILL
XFILL_6_AOI21X1_38 gnd vdd FILL
XFILL_6_AOI21X1_49 gnd vdd FILL
XFILL_73_DFFSR_153 gnd vdd FILL
XFILL_73_DFFSR_164 gnd vdd FILL
XFILL_73_DFFSR_175 gnd vdd FILL
XFILL_16_OAI22X1_18 gnd vdd FILL
XFILL_73_DFFSR_186 gnd vdd FILL
XFILL_6_2 gnd vdd FILL
XFILL_16_OAI22X1_29 gnd vdd FILL
XFILL_73_DFFSR_197 gnd vdd FILL
XFILL_9_NOR2X1_104 gnd vdd FILL
XFILL_77_DFFSR_130 gnd vdd FILL
XFILL_9_NOR2X1_115 gnd vdd FILL
XFILL_9_NOR2X1_126 gnd vdd FILL
XFILL_77_DFFSR_141 gnd vdd FILL
XFILL_77_DFFSR_152 gnd vdd FILL
XFILL_62_4 gnd vdd FILL
XFILL_9_NOR2X1_137 gnd vdd FILL
XFILL_9_NOR2X1_148 gnd vdd FILL
XFILL_77_DFFSR_163 gnd vdd FILL
XFILL_0_CLKBUF1_19 gnd vdd FILL
XFILL_9_NOR2X1_159 gnd vdd FILL
XFILL_77_DFFSR_174 gnd vdd FILL
XFILL_15_NAND3X1_50 gnd vdd FILL
XFILL_77_DFFSR_185 gnd vdd FILL
XFILL_15_NAND3X1_61 gnd vdd FILL
XFILL_77_DFFSR_196 gnd vdd FILL
XFILL_15_NAND3X1_72 gnd vdd FILL
XFILL_28_DFFSR_209 gnd vdd FILL
XFILL_14_AND2X2_3 gnd vdd FILL
XFILL_15_NAND3X1_83 gnd vdd FILL
XFILL_15_NAND3X1_94 gnd vdd FILL
XFILL_36_5_2 gnd vdd FILL
XFILL_35_0_1 gnd vdd FILL
XFILL_1_NAND2X1_2 gnd vdd FILL
XFILL_55_DFFSR_109 gnd vdd FILL
XFILL_11_BUFX4_20 gnd vdd FILL
XFILL_11_BUFX4_31 gnd vdd FILL
XFILL_11_BUFX4_42 gnd vdd FILL
XFILL_5_NAND2X1_1 gnd vdd FILL
XFILL_59_DFFSR_108 gnd vdd FILL
XFILL_11_BUFX4_53 gnd vdd FILL
XFILL_11_BUFX4_64 gnd vdd FILL
XFILL_59_DFFSR_119 gnd vdd FILL
XFILL_11_BUFX4_75 gnd vdd FILL
XFILL_11_BUFX4_86 gnd vdd FILL
XFILL_6_OAI22X1_13 gnd vdd FILL
XFILL_11_BUFX4_97 gnd vdd FILL
XFILL_6_OAI22X1_24 gnd vdd FILL
XFILL_6_OAI22X1_35 gnd vdd FILL
XDFFSR_12 INVX1_32/A DFFSR_7/CLK DFFSR_25/R vdd DFFSR_12/D gnd vdd DFFSR
XFILL_6_OAI22X1_46 gnd vdd FILL
XDFFSR_23 INVX1_28/A DFFSR_4/CLK DFFSR_23/R vdd DFFSR_23/D gnd vdd DFFSR
XFILL_14_NAND3X1_130 gnd vdd FILL
XDFFSR_34 INVX1_27/A CLKBUF1_5/Y DFFSR_49/R vdd DFFSR_34/D gnd vdd DFFSR
XDFFSR_45 INVX1_12/A DFFSR_45/CLK DFFSR_45/R vdd DFFSR_45/D gnd vdd DFFSR
XDFFSR_56 INVX1_5/A DFFSR_56/CLK DFFSR_56/R vdd DFFSR_56/D gnd vdd DFFSR
XFILL_13_DFFSR_220 gnd vdd FILL
XDFFSR_67 DFFSR_67/Q DFFSR_72/CLK DFFSR_96/R vdd DFFSR_67/D gnd vdd DFFSR
XFILL_13_DFFSR_231 gnd vdd FILL
XDFFSR_78 DFFSR_78/Q DFFSR_78/CLK DFFSR_78/R vdd DFFSR_78/D gnd vdd DFFSR
XFILL_13_DFFSR_242 gnd vdd FILL
XDFFSR_89 DFFSR_89/Q CLKBUF1_1/Y DFFSR_89/R vdd DFFSR_89/D gnd vdd DFFSR
XFILL_13_DFFSR_253 gnd vdd FILL
XFILL_13_DFFSR_264 gnd vdd FILL
XFILL_13_DFFSR_275 gnd vdd FILL
XFILL_3_NOR2X1_204 gnd vdd FILL
XFILL_40_DFFSR_120 gnd vdd FILL
XFILL_40_DFFSR_131 gnd vdd FILL
XFILL_1_AOI21X1_7 gnd vdd FILL
XFILL_17_DFFSR_230 gnd vdd FILL
XFILL_5_INVX1_10 gnd vdd FILL
XFILL_40_DFFSR_142 gnd vdd FILL
XFILL_9_NAND2X1_80 gnd vdd FILL
XFILL_5_INVX1_21 gnd vdd FILL
XFILL_5_NAND3X1_102 gnd vdd FILL
XFILL_17_DFFSR_241 gnd vdd FILL
XCLKBUF1_10 BUFX4_84/Y gnd DFFSR_94/CLK vdd CLKBUF1
XFILL_14_BUFX4_9 gnd vdd FILL
XFILL_40_DFFSR_153 gnd vdd FILL
XFILL_5_INVX1_32 gnd vdd FILL
XFILL_9_NAND2X1_91 gnd vdd FILL
XFILL_17_DFFSR_252 gnd vdd FILL
XCLKBUF1_21 BUFX4_9/Y gnd DFFSR_90/CLK vdd CLKBUF1
XFILL_5_NAND3X1_113 gnd vdd FILL
XFILL_5_INVX1_43 gnd vdd FILL
XFILL_17_DFFSR_263 gnd vdd FILL
XFILL_40_DFFSR_164 gnd vdd FILL
XCLKBUF1_32 BUFX4_4/Y gnd DFFSR_7/CLK vdd CLKBUF1
XFILL_40_DFFSR_175 gnd vdd FILL
XFILL_5_NAND3X1_124 gnd vdd FILL
XFILL_5_INVX1_54 gnd vdd FILL
XFILL_6_AND2X2_2 gnd vdd FILL
XFILL_17_DFFSR_274 gnd vdd FILL
XFILL_40_DFFSR_186 gnd vdd FILL
XFILL_5_INVX1_65 gnd vdd FILL
XFILL_14_MUX2X1_19 gnd vdd FILL
XFILL_17_CLKBUF1_11 gnd vdd FILL
XFILL_40_DFFSR_197 gnd vdd FILL
XFILL_5_INVX1_76 gnd vdd FILL
XFILL_17_CLKBUF1_22 gnd vdd FILL
XFILL_5_INVX1_87 gnd vdd FILL
XFILL_44_DFFSR_130 gnd vdd FILL
XFILL_5_INVX1_98 gnd vdd FILL
XFILL_5_AOI21X1_6 gnd vdd FILL
XFILL_17_CLKBUF1_33 gnd vdd FILL
XFILL_44_DFFSR_141 gnd vdd FILL
XFILL_44_DFFSR_152 gnd vdd FILL
XFILL_12_AOI21X1_30 gnd vdd FILL
XFILL_44_DFFSR_163 gnd vdd FILL
XFILL_44_DFFSR_174 gnd vdd FILL
XFILL_12_MUX2X1_8 gnd vdd FILL
XFILL_12_AOI21X1_41 gnd vdd FILL
XFILL_2_DFFSR_1 gnd vdd FILL
XFILL_44_DFFSR_185 gnd vdd FILL
XFILL_27_5_2 gnd vdd FILL
XFILL_18_MUX2X1_18 gnd vdd FILL
XFILL_12_AOI21X1_52 gnd vdd FILL
XFILL_2_5_2 gnd vdd FILL
XFILL_44_DFFSR_196 gnd vdd FILL
XFILL_18_MUX2X1_29 gnd vdd FILL
XFILL_12_AOI21X1_63 gnd vdd FILL
XFILL_12_AOI21X1_74 gnd vdd FILL
XFILL_26_0_1 gnd vdd FILL
XFILL_9_AOI21X1_5 gnd vdd FILL
XFILL_1_0_1 gnd vdd FILL
XFILL_48_DFFSR_140 gnd vdd FILL
XFILL_3_BUFX4_30 gnd vdd FILL
XFILL_3_BUFX4_41 gnd vdd FILL
XFILL_48_DFFSR_151 gnd vdd FILL
XFILL_10_AOI22X1_3 gnd vdd FILL
XFILL_48_DFFSR_162 gnd vdd FILL
XFILL_3_BUFX4_52 gnd vdd FILL
XFILL_3_BUFX4_63 gnd vdd FILL
XFILL_48_DFFSR_173 gnd vdd FILL
XFILL_48_DFFSR_184 gnd vdd FILL
XFILL_3_BUFX4_74 gnd vdd FILL
XFILL_3_BUFX4_85 gnd vdd FILL
XFILL_48_DFFSR_195 gnd vdd FILL
XFILL_22_DFFSR_109 gnd vdd FILL
XFILL_3_BUFX4_96 gnd vdd FILL
XFILL_10_BUFX2_5 gnd vdd FILL
XFILL_14_AOI22X1_2 gnd vdd FILL
XFILL_10_4_2 gnd vdd FILL
XFILL_26_DFFSR_108 gnd vdd FILL
XFILL_26_DFFSR_119 gnd vdd FILL
XFILL_21_MUX2X1_6 gnd vdd FILL
XFILL_18_AOI22X1_1 gnd vdd FILL
XINVX1_106 INVX1_106/A gnd OAI22X1_7/C vdd INVX1
XFILL_0_NAND3X1_120 gnd vdd FILL
XFILL_37_DFFSR_3 gnd vdd FILL
XFILL_0_NAND3X1_131 gnd vdd FILL
XINVX1_117 DFFSR_35/Q gnd NOR3X1_33/A vdd INVX1
XFILL_5_NOR2X1_9 gnd vdd FILL
XINVX1_128 INVX1_128/A gnd INVX1_128/Y vdd INVX1
XINVX1_139 INVX1_139/A gnd INVX1_139/Y vdd INVX1
XFILL_29_DFFSR_10 gnd vdd FILL
XFILL_29_DFFSR_21 gnd vdd FILL
XFILL_15_MUX2X1_102 gnd vdd FILL
XFILL_29_DFFSR_32 gnd vdd FILL
XFILL_29_DFFSR_43 gnd vdd FILL
XFILL_15_MUX2X1_113 gnd vdd FILL
XFILL_15_MUX2X1_124 gnd vdd FILL
XFILL_29_DFFSR_54 gnd vdd FILL
XFILL_15_MUX2X1_135 gnd vdd FILL
XFILL_15_MUX2X1_146 gnd vdd FILL
XFILL_29_DFFSR_65 gnd vdd FILL
XFILL_29_DFFSR_76 gnd vdd FILL
XFILL_29_DFFSR_87 gnd vdd FILL
XFILL_9_1_1 gnd vdd FILL
XFILL_15_MUX2X1_157 gnd vdd FILL
XFILL_29_DFFSR_98 gnd vdd FILL
XFILL_15_MUX2X1_168 gnd vdd FILL
XFILL_2_AOI21X1_80 gnd vdd FILL
XFILL_15_MUX2X1_179 gnd vdd FILL
XFILL_69_DFFSR_20 gnd vdd FILL
XFILL_69_DFFSR_31 gnd vdd FILL
XFILL_72_DFFSR_209 gnd vdd FILL
XFILL_69_DFFSR_42 gnd vdd FILL
XFILL_4_MUX2X1_7 gnd vdd FILL
XFILL_69_DFFSR_53 gnd vdd FILL
XFILL_69_DFFSR_64 gnd vdd FILL
XFILL_69_DFFSR_75 gnd vdd FILL
XFILL_21_DFFSR_9 gnd vdd FILL
XFILL_69_DFFSR_86 gnd vdd FILL
XFILL_26_NOR3X1_19 gnd vdd FILL
XFILL_69_DFFSR_97 gnd vdd FILL
XFILL_5_NOR2X1_190 gnd vdd FILL
XFILL_76_DFFSR_208 gnd vdd FILL
XFILL_11_DFFSR_130 gnd vdd FILL
XFILL_76_DFFSR_219 gnd vdd FILL
XFILL_18_5_2 gnd vdd FILL
XFILL_59_DFFSR_7 gnd vdd FILL
XFILL_11_DFFSR_141 gnd vdd FILL
XFILL_11_DFFSR_152 gnd vdd FILL
XFILL_38_DFFSR_30 gnd vdd FILL
XFILL_11_DFFSR_163 gnd vdd FILL
XFILL_17_0_1 gnd vdd FILL
XFILL_11_DFFSR_174 gnd vdd FILL
XFILL_38_DFFSR_41 gnd vdd FILL
XFILL_0_CLKBUF1_6 gnd vdd FILL
XFILL_38_DFFSR_52 gnd vdd FILL
XFILL_11_DFFSR_185 gnd vdd FILL
XFILL_38_DFFSR_63 gnd vdd FILL
XFILL_38_DFFSR_74 gnd vdd FILL
XFILL_11_DFFSR_196 gnd vdd FILL
XFILL_38_DFFSR_85 gnd vdd FILL
XFILL_15_DFFSR_140 gnd vdd FILL
XFILL_38_DFFSR_96 gnd vdd FILL
XFILL_60_3_2 gnd vdd FILL
XFILL_15_DFFSR_151 gnd vdd FILL
XFILL_27_7 gnd vdd FILL
XFILL_15_DFFSR_162 gnd vdd FILL
XFILL_78_DFFSR_40 gnd vdd FILL
XFILL_15_DFFSR_173 gnd vdd FILL
XFILL_4_CLKBUF1_5 gnd vdd FILL
XFILL_15_DFFSR_184 gnd vdd FILL
XFILL_78_DFFSR_51 gnd vdd FILL
XFILL_22_MUX2X1_170 gnd vdd FILL
XFILL_78_DFFSR_62 gnd vdd FILL
XFILL_15_DFFSR_195 gnd vdd FILL
XFILL_78_DFFSR_73 gnd vdd FILL
XFILL_22_MUX2X1_181 gnd vdd FILL
XFILL_78_DFFSR_84 gnd vdd FILL
XFILL_22_MUX2X1_192 gnd vdd FILL
XFILL_5_MUX2X1_130 gnd vdd FILL
XFILL_78_DFFSR_95 gnd vdd FILL
XFILL_5_MUX2X1_141 gnd vdd FILL
XFILL_19_DFFSR_150 gnd vdd FILL
XFILL_5_MUX2X1_152 gnd vdd FILL
XFILL_5_MUX2X1_163 gnd vdd FILL
XFILL_0_BUFX4_100 gnd vdd FILL
XFILL_19_DFFSR_161 gnd vdd FILL
XFILL_5_MUX2X1_174 gnd vdd FILL
XFILL_19_DFFSR_172 gnd vdd FILL
XFILL_8_CLKBUF1_4 gnd vdd FILL
XFILL_5_MUX2X1_185 gnd vdd FILL
XFILL_19_DFFSR_183 gnd vdd FILL
XFILL_1_INVX1_80 gnd vdd FILL
XFILL_19_DFFSR_194 gnd vdd FILL
XFILL_1_INVX1_91 gnd vdd FILL
XFILL_11_NOR3X1_30 gnd vdd FILL
XFILL_18_NOR3X1_3 gnd vdd FILL
XFILL_11_NOR3X1_41 gnd vdd FILL
XFILL_11_NOR3X1_52 gnd vdd FILL
XFILL_47_DFFSR_50 gnd vdd FILL
XFILL_47_DFFSR_61 gnd vdd FILL
XFILL_61_DFFSR_230 gnd vdd FILL
XFILL_47_DFFSR_72 gnd vdd FILL
XFILL_47_DFFSR_83 gnd vdd FILL
XFILL_61_DFFSR_241 gnd vdd FILL
XFILL_47_DFFSR_94 gnd vdd FILL
XFILL_61_DFFSR_252 gnd vdd FILL
XFILL_61_DFFSR_263 gnd vdd FILL
XFILL_61_DFFSR_274 gnd vdd FILL
XFILL_15_NOR3X1_40 gnd vdd FILL
XFILL_15_NOR3X1_51 gnd vdd FILL
XFILL_87_DFFSR_60 gnd vdd FILL
XFILL_87_DFFSR_71 gnd vdd FILL
XFILL_87_DFFSR_82 gnd vdd FILL
XFILL_65_DFFSR_240 gnd vdd FILL
XFILL_87_DFFSR_93 gnd vdd FILL
XFILL_65_DFFSR_251 gnd vdd FILL
XFILL_65_DFFSR_262 gnd vdd FILL
XFILL_20_CLKBUF1_3 gnd vdd FILL
XFILL_65_DFFSR_273 gnd vdd FILL
XFILL_16_DFFSR_60 gnd vdd FILL
XFILL_11_NAND2X1_18 gnd vdd FILL
XFILL_16_DFFSR_71 gnd vdd FILL
XFILL_16_DFFSR_82 gnd vdd FILL
XFILL_11_NAND2X1_29 gnd vdd FILL
XFILL_19_NOR3X1_50 gnd vdd FILL
XFILL_16_DFFSR_93 gnd vdd FILL
XFILL_60_1 gnd vdd FILL
XFILL_27_NOR3X1_1 gnd vdd FILL
XFILL_69_DFFSR_250 gnd vdd FILL
XFILL_69_DFFSR_261 gnd vdd FILL
XFILL_69_DFFSR_272 gnd vdd FILL
XFILL_24_CLKBUF1_2 gnd vdd FILL
XFILL_56_DFFSR_70 gnd vdd FILL
XFILL_56_DFFSR_81 gnd vdd FILL
XFILL_56_DFFSR_92 gnd vdd FILL
XFILL_43_DFFSR_208 gnd vdd FILL
XFILL_2_NOR2X1_12 gnd vdd FILL
XFILL_8_NAND3X1_11 gnd vdd FILL
XFILL_2_NOR2X1_23 gnd vdd FILL
XFILL_8_NAND3X1_22 gnd vdd FILL
XFILL_43_DFFSR_219 gnd vdd FILL
XFILL_5_OAI21X1_9 gnd vdd FILL
XFILL_2_NOR2X1_34 gnd vdd FILL
XFILL_8_NAND3X1_33 gnd vdd FILL
XFILL_2_NOR2X1_45 gnd vdd FILL
XFILL_1_NOR2X1_2 gnd vdd FILL
XFILL_8_NAND3X1_44 gnd vdd FILL
XFILL_2_NOR2X1_56 gnd vdd FILL
XFILL_8_NAND3X1_55 gnd vdd FILL
XFILL_2_NOR2X1_67 gnd vdd FILL
XFILL_8_NAND3X1_66 gnd vdd FILL
XFILL_2_NOR2X1_78 gnd vdd FILL
XFILL_28_CLKBUF1_1 gnd vdd FILL
XFILL_8_NAND3X1_77 gnd vdd FILL
XFILL_51_3_2 gnd vdd FILL
XFILL_2_NOR2X1_89 gnd vdd FILL
XFILL_8_NAND3X1_88 gnd vdd FILL
XFILL_6_NOR2X1_11 gnd vdd FILL
XFILL_47_DFFSR_207 gnd vdd FILL
XFILL_70_DFFSR_108 gnd vdd FILL
XFILL_8_NAND3X1_99 gnd vdd FILL
XFILL_70_DFFSR_119 gnd vdd FILL
XFILL_47_DFFSR_218 gnd vdd FILL
XFILL_6_NOR2X1_22 gnd vdd FILL
XFILL_9_OAI21X1_8 gnd vdd FILL
XFILL_6_NOR2X1_33 gnd vdd FILL
XFILL_6_NOR2X1_44 gnd vdd FILL
XFILL_47_DFFSR_229 gnd vdd FILL
XFILL_25_DFFSR_80 gnd vdd FILL
XFILL_6_NOR2X1_55 gnd vdd FILL
XFILL_10_OAI22X1_6 gnd vdd FILL
XFILL_25_DFFSR_91 gnd vdd FILL
XFILL_6_NOR2X1_66 gnd vdd FILL
XFILL_6_NOR2X1_77 gnd vdd FILL
XFILL_20_7_0 gnd vdd FILL
XFILL_6_NOR2X1_88 gnd vdd FILL
XFILL_6_NOR2X1_99 gnd vdd FILL
XFILL_74_DFFSR_107 gnd vdd FILL
XFILL_74_DFFSR_118 gnd vdd FILL
XFILL_74_DFFSR_129 gnd vdd FILL
XFILL_14_OAI22X1_5 gnd vdd FILL
XFILL_15_AOI21X1_18 gnd vdd FILL
XFILL_65_DFFSR_90 gnd vdd FILL
XFILL_1_NAND2X1_13 gnd vdd FILL
XFILL_15_AOI21X1_29 gnd vdd FILL
XFILL_15_NAND3X1_120 gnd vdd FILL
XFILL_1_NAND2X1_24 gnd vdd FILL
XFILL_6_DFFSR_2 gnd vdd FILL
XFILL_1_NAND2X1_35 gnd vdd FILL
XFILL_78_DFFSR_106 gnd vdd FILL
XFILL_15_NAND3X1_131 gnd vdd FILL
XFILL_1_NAND2X1_46 gnd vdd FILL
XFILL_1_NAND2X1_57 gnd vdd FILL
XFILL_78_DFFSR_117 gnd vdd FILL
XFILL_76_DFFSR_1 gnd vdd FILL
XFILL_1_NAND2X1_68 gnd vdd FILL
XFILL_78_DFFSR_128 gnd vdd FILL
XFILL_1_NAND2X1_79 gnd vdd FILL
XFILL_78_DFFSR_139 gnd vdd FILL
XFILL_18_OAI22X1_4 gnd vdd FILL
XFILL_8_DFFSR_70 gnd vdd FILL
XFILL_8_DFFSR_81 gnd vdd FILL
XFILL_8_DFFSR_92 gnd vdd FILL
XFILL_1_BUFX2_8 gnd vdd FILL
XFILL_59_4_2 gnd vdd FILL
XFILL_6_NAND3X1_103 gnd vdd FILL
XFILL_32_DFFSR_240 gnd vdd FILL
XFILL_32_DFFSR_251 gnd vdd FILL
XFILL_6_NAND3X1_114 gnd vdd FILL
XFILL_32_DFFSR_262 gnd vdd FILL
XFILL_6_NAND3X1_125 gnd vdd FILL
XFILL_32_DFFSR_273 gnd vdd FILL
XFILL_27_CLKBUF1_12 gnd vdd FILL
XFILL_27_CLKBUF1_23 gnd vdd FILL
XFILL_27_CLKBUF1_34 gnd vdd FILL
XFILL_60_DFFSR_7 gnd vdd FILL
XFILL_36_DFFSR_250 gnd vdd FILL
XFILL_1_AOI22X1_11 gnd vdd FILL
XFILL_36_DFFSR_261 gnd vdd FILL
XFILL_36_DFFSR_272 gnd vdd FILL
XFILL_2_MUX2X1_30 gnd vdd FILL
XFILL_2_MUX2X1_41 gnd vdd FILL
XFILL_10_DFFSR_208 gnd vdd FILL
XFILL_5_AOI21X1_13 gnd vdd FILL
XFILL_2_MUX2X1_52 gnd vdd FILL
XFILL_10_DFFSR_219 gnd vdd FILL
XFILL_42_3_2 gnd vdd FILL
XFILL_5_AOI21X1_24 gnd vdd FILL
XFILL_2_MUX2X1_63 gnd vdd FILL
XFILL_63_DFFSR_150 gnd vdd FILL
XFILL_2_MUX2X1_74 gnd vdd FILL
XFILL_5_AOI21X1_35 gnd vdd FILL
XFILL_5_AOI21X1_46 gnd vdd FILL
XFILL_2_MUX2X1_85 gnd vdd FILL
XFILL_63_DFFSR_161 gnd vdd FILL
XFILL_2_MUX2X1_96 gnd vdd FILL
XFILL_5_AOI21X1_57 gnd vdd FILL
XFILL_5_AOI21X1_68 gnd vdd FILL
XFILL_63_DFFSR_172 gnd vdd FILL
XFILL_15_OAI22X1_15 gnd vdd FILL
XFILL_63_DFFSR_183 gnd vdd FILL
XFILL_15_OAI22X1_26 gnd vdd FILL
XFILL_63_DFFSR_194 gnd vdd FILL
XFILL_5_AOI21X1_79 gnd vdd FILL
XFILL_15_OAI22X1_37 gnd vdd FILL
XFILL_14_DFFSR_207 gnd vdd FILL
XFILL_6_MUX2X1_40 gnd vdd FILL
XFILL_8_NOR2X1_101 gnd vdd FILL
XFILL_15_OAI22X1_48 gnd vdd FILL
XFILL_6_MUX2X1_51 gnd vdd FILL
XFILL_11_NAND3X1_7 gnd vdd FILL
XFILL_6_MUX2X1_62 gnd vdd FILL
XFILL_11_7_0 gnd vdd FILL
XFILL_14_DFFSR_218 gnd vdd FILL
XFILL_8_NOR2X1_112 gnd vdd FILL
XFILL_8_NOR2X1_123 gnd vdd FILL
XFILL_14_DFFSR_229 gnd vdd FILL
XFILL_6_MUX2X1_73 gnd vdd FILL
XFILL_8_NOR2X1_134 gnd vdd FILL
XFILL_0_BUFX4_2 gnd vdd FILL
XFILL_67_DFFSR_160 gnd vdd FILL
XFILL_8_NOR2X1_145 gnd vdd FILL
XFILL_6_MUX2X1_84 gnd vdd FILL
XFILL_6_MUX2X1_95 gnd vdd FILL
XFILL_8_NOR2X1_156 gnd vdd FILL
XFILL_4_BUFX4_19 gnd vdd FILL
XFILL_67_DFFSR_171 gnd vdd FILL
XFILL_8_NOR2X1_167 gnd vdd FILL
XFILL_67_DFFSR_182 gnd vdd FILL
XFILL_8_NOR2X1_178 gnd vdd FILL
XFILL_67_DFFSR_193 gnd vdd FILL
XFILL_18_DFFSR_206 gnd vdd FILL
XFILL_41_DFFSR_107 gnd vdd FILL
XFILL_8_NOR2X1_189 gnd vdd FILL
XFILL_18_DFFSR_217 gnd vdd FILL
XFILL_41_DFFSR_118 gnd vdd FILL
XFILL_15_NAND3X1_6 gnd vdd FILL
XFILL_14_NAND3X1_80 gnd vdd FILL
XFILL_41_DFFSR_129 gnd vdd FILL
XFILL_14_NAND3X1_91 gnd vdd FILL
XFILL_18_DFFSR_228 gnd vdd FILL
XFILL_18_DFFSR_239 gnd vdd FILL
XFILL_1_NAND3X1_110 gnd vdd FILL
XFILL_1_NAND3X1_121 gnd vdd FILL
XFILL_1_NAND3X1_132 gnd vdd FILL
XFILL_45_DFFSR_106 gnd vdd FILL
XFILL_45_DFFSR_117 gnd vdd FILL
XFILL_45_DFFSR_128 gnd vdd FILL
XFILL_45_DFFSR_139 gnd vdd FILL
XFILL_49_DFFSR_105 gnd vdd FILL
XFILL_8_MUX2X1_107 gnd vdd FILL
XFILL_8_MUX2X1_118 gnd vdd FILL
XFILL_49_DFFSR_116 gnd vdd FILL
XFILL_8_MUX2X1_129 gnd vdd FILL
XFILL_49_DFFSR_127 gnd vdd FILL
XFILL_49_DFFSR_138 gnd vdd FILL
XFILL_49_DFFSR_149 gnd vdd FILL
XFILL_5_OAI22X1_10 gnd vdd FILL
XFILL_11_AND2X2_7 gnd vdd FILL
XFILL_22_MUX2X1_60 gnd vdd FILL
XFILL_5_OAI22X1_21 gnd vdd FILL
XFILL_22_MUX2X1_71 gnd vdd FILL
XFILL_22_MUX2X1_82 gnd vdd FILL
XFILL_5_OAI22X1_32 gnd vdd FILL
XFILL_5_OAI22X1_43 gnd vdd FILL
XFILL_22_MUX2X1_93 gnd vdd FILL
XFILL_9_OAI21X1_12 gnd vdd FILL
XFILL_9_OAI21X1_23 gnd vdd FILL
XFILL_9_OAI21X1_34 gnd vdd FILL
XFILL_9_OAI21X1_45 gnd vdd FILL
XFILL_32_5 gnd vdd FILL
XFILL_61_6_0 gnd vdd FILL
XFILL_33_3_2 gnd vdd FILL
XFILL_2_NOR2X1_201 gnd vdd FILL
XFILL_25_4 gnd vdd FILL
XFILL_30_DFFSR_150 gnd vdd FILL
XFILL_18_3 gnd vdd FILL
XFILL_30_DFFSR_161 gnd vdd FILL
XFILL_30_DFFSR_172 gnd vdd FILL
XFILL_30_DFFSR_183 gnd vdd FILL
XFILL_30_DFFSR_194 gnd vdd FILL
XFILL_39_DFFSR_19 gnd vdd FILL
XFILL_16_CLKBUF1_30 gnd vdd FILL
XFILL_16_CLKBUF1_41 gnd vdd FILL
XFILL_34_DFFSR_160 gnd vdd FILL
XFILL_34_DFFSR_171 gnd vdd FILL
XFILL_34_DFFSR_182 gnd vdd FILL
XFILL_34_DFFSR_193 gnd vdd FILL
XFILL_79_DFFSR_18 gnd vdd FILL
XFILL_11_AOI21X1_60 gnd vdd FILL
XFILL_11_AOI21X1_71 gnd vdd FILL
XFILL_79_DFFSR_29 gnd vdd FILL
XFILL_38_DFFSR_170 gnd vdd FILL
XFILL_2_INVX1_14 gnd vdd FILL
XFILL_2_INVX1_25 gnd vdd FILL
XFILL_38_DFFSR_181 gnd vdd FILL
XFILL_2_INVX1_36 gnd vdd FILL
XFILL_38_DFFSR_192 gnd vdd FILL
XFILL_12_DFFSR_106 gnd vdd FILL
XFILL_2_INVX1_47 gnd vdd FILL
XFILL_12_DFFSR_117 gnd vdd FILL
XFILL_2_INVX1_58 gnd vdd FILL
XFILL_3_AND2X2_6 gnd vdd FILL
XFILL_30_NOR3X1_50 gnd vdd FILL
XFILL_12_DFFSR_128 gnd vdd FILL
XFILL_2_INVX1_69 gnd vdd FILL
XFILL_12_DFFSR_139 gnd vdd FILL
XFILL_48_DFFSR_17 gnd vdd FILL
XFILL_48_DFFSR_28 gnd vdd FILL
XFILL_48_DFFSR_39 gnd vdd FILL
XFILL_80_DFFSR_250 gnd vdd FILL
XFILL_80_DFFSR_261 gnd vdd FILL
XFILL_16_DFFSR_105 gnd vdd FILL
XFILL_80_DFFSR_272 gnd vdd FILL
XFILL_16_DFFSR_116 gnd vdd FILL
XFILL_16_DFFSR_127 gnd vdd FILL
XFILL_16_DFFSR_138 gnd vdd FILL
XFILL_16_DFFSR_149 gnd vdd FILL
XFILL_11_AOI21X1_1 gnd vdd FILL
XFILL_0_BUFX4_12 gnd vdd FILL
XFILL_42_DFFSR_4 gnd vdd FILL
XFILL_0_BUFX4_23 gnd vdd FILL
XFILL_0_BUFX4_34 gnd vdd FILL
XFILL_0_BUFX4_45 gnd vdd FILL
XFILL_84_DFFSR_260 gnd vdd FILL
XFILL_84_DFFSR_271 gnd vdd FILL
XFILL_17_DFFSR_16 gnd vdd FILL
XFILL_17_DFFSR_27 gnd vdd FILL
XFILL_0_BUFX4_56 gnd vdd FILL
XFILL_17_DFFSR_38 gnd vdd FILL
XFILL_0_BUFX4_67 gnd vdd FILL
XFILL_0_BUFX4_78 gnd vdd FILL
XFILL_14_MUX2X1_110 gnd vdd FILL
XFILL_17_DFFSR_49 gnd vdd FILL
XFILL_0_BUFX4_89 gnd vdd FILL
XFILL_14_MUX2X1_121 gnd vdd FILL
XFILL_52_6_0 gnd vdd FILL
XFILL_14_MUX2X1_132 gnd vdd FILL
XFILL_24_3_2 gnd vdd FILL
XFILL_14_MUX2X1_143 gnd vdd FILL
XFILL_14_MUX2X1_154 gnd vdd FILL
XFILL_12_NOR3X1_17 gnd vdd FILL
XFILL_14_MUX2X1_165 gnd vdd FILL
XFILL_57_DFFSR_15 gnd vdd FILL
XFILL_5_BUFX2_9 gnd vdd FILL
XFILL_12_NOR3X1_28 gnd vdd FILL
XFILL_57_DFFSR_26 gnd vdd FILL
XFILL_14_MUX2X1_176 gnd vdd FILL
XFILL_14_MUX2X1_187 gnd vdd FILL
XFILL_57_DFFSR_37 gnd vdd FILL
XFILL_12_NOR3X1_39 gnd vdd FILL
XFILL_62_DFFSR_206 gnd vdd FILL
XFILL_57_DFFSR_48 gnd vdd FILL
XFILL_62_DFFSR_217 gnd vdd FILL
XFILL_57_DFFSR_59 gnd vdd FILL
XFILL_62_DFFSR_228 gnd vdd FILL
XFILL_62_DFFSR_239 gnd vdd FILL
XFILL_16_NOR3X1_16 gnd vdd FILL
XFILL_16_NOR3X1_27 gnd vdd FILL
XFILL_16_NOR3X1_38 gnd vdd FILL
XFILL_16_NOR3X1_49 gnd vdd FILL
XFILL_66_DFFSR_205 gnd vdd FILL
XFILL_64_DFFSR_8 gnd vdd FILL
XFILL_66_DFFSR_216 gnd vdd FILL
XFILL_26_DFFSR_14 gnd vdd FILL
XFILL_66_DFFSR_227 gnd vdd FILL
XFILL_26_DFFSR_25 gnd vdd FILL
XFILL_26_DFFSR_36 gnd vdd FILL
XFILL_66_DFFSR_238 gnd vdd FILL
XFILL_66_DFFSR_249 gnd vdd FILL
XFILL_26_DFFSR_47 gnd vdd FILL
XFILL_26_DFFSR_58 gnd vdd FILL
XFILL_26_DFFSR_69 gnd vdd FILL
XFILL_66_DFFSR_13 gnd vdd FILL
XFILL_66_DFFSR_24 gnd vdd FILL
XFILL_66_DFFSR_35 gnd vdd FILL
XFILL_66_DFFSR_46 gnd vdd FILL
XFILL_66_DFFSR_57 gnd vdd FILL
XFILL_66_DFFSR_68 gnd vdd FILL
XNAND3X1_12 DFFSR_36/Q BUFX4_5/Y NOR2X1_29/Y gnd NAND3X1_16/A vdd NAND3X1
XFILL_66_DFFSR_79 gnd vdd FILL
XNAND3X1_23 DFFSR_102/Q BUFX4_102/Y NOR2X1_37/Y gnd OAI21X1_31/C vdd NAND3X1
XFILL_7_4_2 gnd vdd FILL
XNAND3X1_34 INVX2_4/Y OAI21X1_41/A OAI21X1_48/A gnd NAND3X1_36/C vdd NAND3X1
XNAND3X1_45 OAI21X1_1/A NAND2X1_4/B AND2X2_8/B gnd MUX2X1_7/S vdd NAND3X1
XFILL_4_BUFX4_3 gnd vdd FILL
XNAND3X1_56 OAI21X1_48/A OAI21X1_12/Y AOI22X1_2/C gnd AOI22X1_1/C vdd NAND3X1
XFILL_4_MUX2X1_160 gnd vdd FILL
XFILL_9_DFFSR_15 gnd vdd FILL
XFILL_9_DFFSR_26 gnd vdd FILL
XFILL_4_MUX2X1_171 gnd vdd FILL
XNAND3X1_67 INVX2_3/A OAI21X1_40/Y OAI21X1_39/Y gnd NAND3X1_67/Y vdd NAND3X1
XFILL_7_NAND3X1_104 gnd vdd FILL
XFILL_35_DFFSR_12 gnd vdd FILL
XFILL_9_DFFSR_37 gnd vdd FILL
XFILL_7_NAND3X1_115 gnd vdd FILL
XNAND3X1_78 INVX2_4/Y OAI21X1_35/A OAI21X1_48/A gnd NAND3X1_78/Y vdd NAND3X1
XNAND3X1_89 NOR3X1_9/B NOR3X1_9/A AND2X2_1/B gnd NOR3X1_1/B vdd NAND3X1
XFILL_9_DFFSR_48 gnd vdd FILL
XFILL_4_MUX2X1_182 gnd vdd FILL
XFILL_35_DFFSR_23 gnd vdd FILL
XFILL_7_NAND3X1_126 gnd vdd FILL
XNOR2X1_12 NOR2X1_12/A NOR2X1_12/B gnd NOR2X1_12/Y vdd NOR2X1
XFILL_9_DFFSR_59 gnd vdd FILL
XFILL_4_MUX2X1_193 gnd vdd FILL
XFILL_35_DFFSR_34 gnd vdd FILL
XNOR2X1_23 NOR2X1_68/A OR2X2_1/A gnd NOR2X1_23/Y vdd NOR2X1
XFILL_35_DFFSR_45 gnd vdd FILL
XFILL_35_DFFSR_56 gnd vdd FILL
XNOR2X1_34 NOR3X1_2/C NOR2X1_44/B gnd NOR2X1_34/Y vdd NOR2X1
XFILL_35_DFFSR_67 gnd vdd FILL
XNOR2X1_45 AND2X2_2/A NOR2X1_45/B gnd BUFX4_92/A vdd NOR2X1
XNOR2X1_56 OAI21X1_4/Y OAI22X1_4/Y gnd NOR2X1_56/Y vdd NOR2X1
XFILL_35_DFFSR_78 gnd vdd FILL
XNOR2X1_67 NOR2X1_67/A OAI21X1_9/Y gnd NOR2X1_67/Y vdd NOR2X1
XFILL_35_DFFSR_89 gnd vdd FILL
XNOR2X1_78 NOR2X1_78/A NOR2X1_78/B gnd NOR2X1_78/Y vdd NOR2X1
XFILL_75_DFFSR_11 gnd vdd FILL
XFILL_75_DFFSR_22 gnd vdd FILL
XFILL_51_DFFSR_260 gnd vdd FILL
XNOR2X1_89 NOR2X1_89/A NOR2X1_89/B gnd NOR2X1_89/Y vdd NOR2X1
XFILL_51_DFFSR_271 gnd vdd FILL
XFILL_43_6_0 gnd vdd FILL
XFILL_75_DFFSR_33 gnd vdd FILL
XFILL_15_3_2 gnd vdd FILL
XFILL_18_MUX2X1_1 gnd vdd FILL
XFILL_75_DFFSR_44 gnd vdd FILL
XFILL_75_DFFSR_55 gnd vdd FILL
XFILL_75_DFFSR_66 gnd vdd FILL
XFILL_75_DFFSR_77 gnd vdd FILL
XFILL_75_DFFSR_88 gnd vdd FILL
XFILL_75_DFFSR_99 gnd vdd FILL
XFILL_3_INVX1_7 gnd vdd FILL
XFILL_55_DFFSR_270 gnd vdd FILL
XFILL_10_NAND2X1_15 gnd vdd FILL
XFILL_10_NAND2X1_26 gnd vdd FILL
XFILL_44_DFFSR_10 gnd vdd FILL
XFILL_10_NAND2X1_37 gnd vdd FILL
XFILL_44_DFFSR_21 gnd vdd FILL
XFILL_10_NAND2X1_48 gnd vdd FILL
XFILL_44_DFFSR_32 gnd vdd FILL
XFILL_44_DFFSR_43 gnd vdd FILL
XFILL_10_NAND2X1_59 gnd vdd FILL
XFILL_15_NOR3X1_7 gnd vdd FILL
XFILL_44_DFFSR_54 gnd vdd FILL
XFILL_44_DFFSR_65 gnd vdd FILL
XFILL_44_DFFSR_76 gnd vdd FILL
XFILL_82_DFFSR_170 gnd vdd FILL
XFILL_44_DFFSR_87 gnd vdd FILL
XFILL_82_DFFSR_181 gnd vdd FILL
XFILL_44_DFFSR_98 gnd vdd FILL
XFILL_82_DFFSR_192 gnd vdd FILL
XFILL_33_DFFSR_205 gnd vdd FILL
XFILL_33_DFFSR_216 gnd vdd FILL
XFILL_84_DFFSR_20 gnd vdd FILL
XFILL_84_DFFSR_31 gnd vdd FILL
XFILL_33_DFFSR_227 gnd vdd FILL
XFILL_84_DFFSR_42 gnd vdd FILL
XFILL_7_NAND3X1_30 gnd vdd FILL
XFILL_2_DFFSR_240 gnd vdd FILL
XFILL_2_NAND3X1_100 gnd vdd FILL
XFILL_2_DFFSR_251 gnd vdd FILL
XFILL_33_DFFSR_238 gnd vdd FILL
XFILL_84_DFFSR_53 gnd vdd FILL
XFILL_7_NAND3X1_41 gnd vdd FILL
XFILL_2_NAND3X1_111 gnd vdd FILL
XFILL_33_DFFSR_249 gnd vdd FILL
XFILL_2_DFFSR_262 gnd vdd FILL
XFILL_13_DFFSR_20 gnd vdd FILL
XFILL_2_DFFSR_273 gnd vdd FILL
XFILL_84_DFFSR_64 gnd vdd FILL
XFILL_2_NAND3X1_122 gnd vdd FILL
XFILL_7_NAND3X1_52 gnd vdd FILL
XFILL_13_DFFSR_31 gnd vdd FILL
XFILL_84_DFFSR_75 gnd vdd FILL
XFILL_7_NAND3X1_63 gnd vdd FILL
XFILL_86_DFFSR_180 gnd vdd FILL
XFILL_84_DFFSR_86 gnd vdd FILL
XFILL_7_NAND3X1_74 gnd vdd FILL
XFILL_13_DFFSR_42 gnd vdd FILL
XFILL_7_NAND3X1_85 gnd vdd FILL
XFILL_13_DFFSR_53 gnd vdd FILL
XFILL_86_DFFSR_191 gnd vdd FILL
XFILL_84_DFFSR_97 gnd vdd FILL
XFILL_7_NAND3X1_96 gnd vdd FILL
XFILL_60_DFFSR_105 gnd vdd FILL
XFILL_37_DFFSR_204 gnd vdd FILL
XFILL_37_DFFSR_215 gnd vdd FILL
XFILL_60_DFFSR_116 gnd vdd FILL
XFILL_13_DFFSR_64 gnd vdd FILL
XFILL_60_DFFSR_127 gnd vdd FILL
XFILL_37_DFFSR_226 gnd vdd FILL
XFILL_13_DFFSR_75 gnd vdd FILL
XFILL_60_DFFSR_138 gnd vdd FILL
XFILL_13_DFFSR_86 gnd vdd FILL
XFILL_7_INVX8_1 gnd vdd FILL
XFILL_37_DFFSR_237 gnd vdd FILL
XFILL_6_DFFSR_250 gnd vdd FILL
XFILL_13_DFFSR_97 gnd vdd FILL
XFILL_60_DFFSR_149 gnd vdd FILL
XFILL_37_DFFSR_248 gnd vdd FILL
XFILL_6_DFFSR_261 gnd vdd FILL
XFILL_6_DFFSR_272 gnd vdd FILL
XFILL_37_DFFSR_259 gnd vdd FILL
XFILL_53_DFFSR_30 gnd vdd FILL
XFILL_53_DFFSR_41 gnd vdd FILL
XFILL_3_MUX2X1_17 gnd vdd FILL
XFILL_24_NOR3X1_5 gnd vdd FILL
XFILL_64_DFFSR_104 gnd vdd FILL
XFILL_53_DFFSR_52 gnd vdd FILL
XFILL_3_MUX2X1_28 gnd vdd FILL
XFILL_53_DFFSR_63 gnd vdd FILL
XFILL_3_MUX2X1_39 gnd vdd FILL
XFILL_19_CLKBUF1_18 gnd vdd FILL
XFILL_64_DFFSR_115 gnd vdd FILL
XFILL_19_CLKBUF1_29 gnd vdd FILL
XFILL_53_DFFSR_74 gnd vdd FILL
XFILL_64_DFFSR_126 gnd vdd FILL
XFILL_64_DFFSR_137 gnd vdd FILL
XFILL_53_DFFSR_85 gnd vdd FILL
XFILL_64_DFFSR_148 gnd vdd FILL
XFILL_53_DFFSR_96 gnd vdd FILL
XFILL_65_2_2 gnd vdd FILL
XFILL_0_NAND2X1_10 gnd vdd FILL
XFILL_14_AOI21X1_15 gnd vdd FILL
XFILL_14_AOI21X1_26 gnd vdd FILL
XFILL_64_DFFSR_159 gnd vdd FILL
XFILL_0_NAND2X1_21 gnd vdd FILL
XFILL_14_AOI21X1_37 gnd vdd FILL
XNOR2X1_102 INVX1_33/Y NOR2X1_51/B gnd NOR2X1_102/Y vdd NOR2X1
XMUX2X1_30 BUFX4_63/Y INVX1_43/Y NOR2X1_19/B gnd MUX2X1_30/Y vdd MUX2X1
XFILL_0_NAND2X1_32 gnd vdd FILL
XFILL_7_MUX2X1_16 gnd vdd FILL
XFILL_14_AOI21X1_48 gnd vdd FILL
XFILL_24_DFFSR_1 gnd vdd FILL
XFILL_68_DFFSR_103 gnd vdd FILL
XMUX2X1_41 INVX1_54/Y MUX2X1_4/B NAND2X1_6/Y gnd MUX2X1_41/Y vdd MUX2X1
XFILL_7_MUX2X1_27 gnd vdd FILL
XFILL_0_NAND2X1_43 gnd vdd FILL
XNOR2X1_113 DFFSR_160/Q NOR2X1_90/B gnd NOR2X1_113/Y vdd NOR2X1
XFILL_14_AOI21X1_59 gnd vdd FILL
XMUX2X1_52 INVX1_65/Y MUX2X1_6/B NAND2X1_8/Y gnd MUX2X1_52/Y vdd MUX2X1
XFILL_7_MUX2X1_38 gnd vdd FILL
XFILL_0_NAND2X1_54 gnd vdd FILL
XNOR2X1_124 DFFSR_148/Q AOI21X1_3/B gnd NOR2X1_124/Y vdd NOR2X1
XFILL_0_NAND2X1_65 gnd vdd FILL
XFILL_68_DFFSR_114 gnd vdd FILL
XMUX2X1_63 BUFX4_85/Y INVX1_76/Y NOR2X1_23/Y gnd MUX2X1_63/Y vdd MUX2X1
XFILL_7_MUX2X1_49 gnd vdd FILL
XFILL_81_DFFSR_2 gnd vdd FILL
XMUX2X1_74 INVX1_87/Y BUFX4_75/Y OR2X2_1/Y gnd MUX2X1_74/Y vdd MUX2X1
XNOR2X1_135 NOR2X1_24/A NOR2X1_138/A gnd INVX1_166/A vdd NOR2X1
XFILL_0_NAND2X1_76 gnd vdd FILL
XFILL_68_DFFSR_125 gnd vdd FILL
XFILL_68_DFFSR_136 gnd vdd FILL
XFILL_22_DFFSR_40 gnd vdd FILL
XNOR2X1_146 NAND3X1_3/A AOI21X1_9/B gnd NOR2X1_146/Y vdd NOR2X1
XFILL_34_6_0 gnd vdd FILL
XFILL_11_OAI21X1_4 gnd vdd FILL
XFILL_22_DFFSR_51 gnd vdd FILL
XMUX2X1_85 INVX1_98/Y BUFX4_75/Y MUX2X1_86/S gnd MUX2X1_85/Y vdd MUX2X1
XFILL_0_NAND2X1_87 gnd vdd FILL
XFILL_68_DFFSR_147 gnd vdd FILL
XFILL_68_DFFSR_158 gnd vdd FILL
XMUX2X1_96 MUX2X1_96/A MUX2X1_8/A MUX2X1_99/S gnd DFFSR_57/D vdd MUX2X1
XNOR2X1_157 NAND2X1_3/Y INVX1_205/Y gnd NOR2X1_161/B vdd NOR2X1
XFILL_22_DFFSR_62 gnd vdd FILL
XFILL_22_DFFSR_73 gnd vdd FILL
XNOR2X1_168 NAND2X1_3/Y INVX1_3/Y gnd NOR2X1_168/Y vdd NOR2X1
XNOR2X1_179 DFFSR_29/Q NOR2X1_181/B gnd NOR2X1_179/Y vdd NOR2X1
XFILL_68_DFFSR_169 gnd vdd FILL
XFILL_22_DFFSR_84 gnd vdd FILL
XFILL_23_1 gnd vdd FILL
XFILL_22_DFFSR_95 gnd vdd FILL
XFILL_7_NOR3X1_6 gnd vdd FILL
XFILL_15_OAI21X1_3 gnd vdd FILL
XFILL_62_DFFSR_50 gnd vdd FILL
XFILL_62_DFFSR_61 gnd vdd FILL
XFILL_62_DFFSR_72 gnd vdd FILL
XFILL_62_DFFSR_83 gnd vdd FILL
XFILL_22_DFFSR_270 gnd vdd FILL
XFILL_62_DFFSR_94 gnd vdd FILL
XFILL_3_INVX1_210 gnd vdd FILL
XFILL_3_INVX1_221 gnd vdd FILL
XFILL_26_CLKBUF1_20 gnd vdd FILL
XFILL_26_CLKBUF1_31 gnd vdd FILL
XFILL_26_CLKBUF1_42 gnd vdd FILL
XFILL_5_DFFSR_30 gnd vdd FILL
XFILL_46_DFFSR_5 gnd vdd FILL
XFILL_5_DFFSR_41 gnd vdd FILL
XFILL_5_DFFSR_52 gnd vdd FILL
XFILL_5_DFFSR_63 gnd vdd FILL
XMUX2X1_108 MUX2X1_2/A INVX1_149/Y NOR2X1_57/Y gnd DFFSR_164/D vdd MUX2X1
XFILL_5_DFFSR_74 gnd vdd FILL
XFILL_9_CLKBUF1_13 gnd vdd FILL
XMUX2X1_119 INVX1_161/Y MUX2X1_1/A NAND2X1_78/Y gnd DFFSR_136/D vdd MUX2X1
XFILL_9_CLKBUF1_24 gnd vdd FILL
XFILL_5_DFFSR_85 gnd vdd FILL
XFILL_31_DFFSR_60 gnd vdd FILL
XFILL_23_MUX2X1_14 gnd vdd FILL
XFILL_7_INVX1_220 gnd vdd FILL
XFILL_23_MUX2X1_25 gnd vdd FILL
XFILL_5_DFFSR_96 gnd vdd FILL
XFILL_9_CLKBUF1_35 gnd vdd FILL
XFILL_31_DFFSR_71 gnd vdd FILL
XFILL_31_DFFSR_82 gnd vdd FILL
XFILL_4_AOI21X1_10 gnd vdd FILL
XFILL_23_MUX2X1_36 gnd vdd FILL
XFILL_17_MUX2X1_109 gnd vdd FILL
XFILL_31_DFFSR_93 gnd vdd FILL
XFILL_4_AOI21X1_21 gnd vdd FILL
XFILL_23_MUX2X1_47 gnd vdd FILL
XFILL_23_MUX2X1_58 gnd vdd FILL
XFILL_4_AOI21X1_32 gnd vdd FILL
XFILL_4_AOI21X1_43 gnd vdd FILL
XFILL_23_MUX2X1_69 gnd vdd FILL
XFILL_4_AOI21X1_54 gnd vdd FILL
XFILL_14_OAI22X1_12 gnd vdd FILL
XFILL_4_AOI21X1_65 gnd vdd FILL
XFILL_53_DFFSR_180 gnd vdd FILL
XFILL_14_OAI22X1_23 gnd vdd FILL
XFILL_4_AOI21X1_76 gnd vdd FILL
XFILL_14_OAI22X1_34 gnd vdd FILL
XFILL_53_DFFSR_191 gnd vdd FILL
XINVX1_15 INVX1_15/A gnd INVX1_15/Y vdd INVX1
XFILL_71_DFFSR_70 gnd vdd FILL
XFILL_14_OAI22X1_45 gnd vdd FILL
XINVX1_26 INVX1_26/A gnd INVX1_26/Y vdd INVX1
XFILL_71_DFFSR_81 gnd vdd FILL
XINVX1_37 INVX1_37/A gnd INVX1_37/Y vdd INVX1
XFILL_71_DFFSR_92 gnd vdd FILL
XFILL_7_NOR2X1_120 gnd vdd FILL
XINVX1_48 INVX1_48/A gnd INVX1_48/Y vdd INVX1
XFILL_7_NOR2X1_131 gnd vdd FILL
XINVX1_59 INVX1_59/A gnd INVX1_59/Y vdd INVX1
XFILL_7_NOR2X1_142 gnd vdd FILL
XFILL_7_NOR2X1_153 gnd vdd FILL
XFILL_7_NOR2X1_164 gnd vdd FILL
XFILL_57_DFFSR_190 gnd vdd FILL
XFILL_7_NOR2X1_175 gnd vdd FILL
XFILL_31_DFFSR_104 gnd vdd FILL
XFILL_56_2_2 gnd vdd FILL
XFILL_7_NOR2X1_186 gnd vdd FILL
XFILL_68_DFFSR_9 gnd vdd FILL
XFILL_7_NOR2X1_197 gnd vdd FILL
XFILL_31_DFFSR_115 gnd vdd FILL
XFILL_31_DFFSR_126 gnd vdd FILL
XFILL_31_DFFSR_137 gnd vdd FILL
XFILL_0_DFFSR_150 gnd vdd FILL
XFILL_31_DFFSR_148 gnd vdd FILL
XFILL_11_NOR2X1_203 gnd vdd FILL
XFILL_0_DFFSR_161 gnd vdd FILL
XFILL_40_DFFSR_80 gnd vdd FILL
XFILL_0_DFFSR_172 gnd vdd FILL
XFILL_31_DFFSR_159 gnd vdd FILL
XFILL_0_DFFSR_183 gnd vdd FILL
XFILL_40_DFFSR_91 gnd vdd FILL
XFILL_0_DFFSR_194 gnd vdd FILL
XFILL_35_DFFSR_103 gnd vdd FILL
XFILL_25_6_0 gnd vdd FILL
XFILL_0_6_0 gnd vdd FILL
XFILL_35_DFFSR_114 gnd vdd FILL
XFILL_35_DFFSR_125 gnd vdd FILL
XFILL_35_DFFSR_136 gnd vdd FILL
XFILL_4_DFFSR_160 gnd vdd FILL
XFILL_35_DFFSR_147 gnd vdd FILL
XFILL_35_DFFSR_158 gnd vdd FILL
XFILL_4_DFFSR_171 gnd vdd FILL
XFILL_80_DFFSR_90 gnd vdd FILL
XFILL_35_DFFSR_169 gnd vdd FILL
XFILL_4_DFFSR_182 gnd vdd FILL
XFILL_4_DFFSR_193 gnd vdd FILL
XFILL_39_DFFSR_102 gnd vdd FILL
XFILL_7_MUX2X1_104 gnd vdd FILL
XFILL_7_MUX2X1_115 gnd vdd FILL
XFILL_39_DFFSR_113 gnd vdd FILL
XFILL_7_MUX2X1_126 gnd vdd FILL
XFILL_39_DFFSR_124 gnd vdd FILL
XFILL_39_DFFSR_135 gnd vdd FILL
XFILL_7_MUX2X1_137 gnd vdd FILL
XFILL_39_DFFSR_146 gnd vdd FILL
XFILL_8_BUFX4_4 gnd vdd FILL
XFILL_7_MUX2X1_148 gnd vdd FILL
XFILL_39_DFFSR_157 gnd vdd FILL
XFILL_8_DFFSR_170 gnd vdd FILL
XFILL_7_MUX2X1_159 gnd vdd FILL
XFILL_39_DFFSR_168 gnd vdd FILL
XFILL_8_DFFSR_181 gnd vdd FILL
XFILL_39_DFFSR_179 gnd vdd FILL
XFILL_12_MUX2X1_90 gnd vdd FILL
XFILL_31_NOR3X1_15 gnd vdd FILL
XFILL_4_OAI22X1_40 gnd vdd FILL
XFILL_8_DFFSR_192 gnd vdd FILL
XFILL_4_OAI22X1_51 gnd vdd FILL
XFILL_31_NOR3X1_26 gnd vdd FILL
XFILL_0_NOR3X1_50 gnd vdd FILL
XFILL_8_OAI21X1_20 gnd vdd FILL
XFILL_31_NOR3X1_37 gnd vdd FILL
XFILL_8_OAI21X1_31 gnd vdd FILL
XFILL_31_NOR3X1_48 gnd vdd FILL
XFILL_81_DFFSR_204 gnd vdd FILL
XFILL_81_DFFSR_215 gnd vdd FILL
XFILL_8_OAI21X1_42 gnd vdd FILL
XFILL_81_DFFSR_226 gnd vdd FILL
XFILL_81_DFFSR_237 gnd vdd FILL
XFILL_81_DFFSR_248 gnd vdd FILL
XFILL_81_DFFSR_259 gnd vdd FILL
XFILL_85_DFFSR_203 gnd vdd FILL
XFILL_85_DFFSR_214 gnd vdd FILL
XFILL_85_DFFSR_225 gnd vdd FILL
XFILL_8_7_0 gnd vdd FILL
XFILL_85_DFFSR_236 gnd vdd FILL
XFILL_7_INVX1_8 gnd vdd FILL
XFILL_85_DFFSR_247 gnd vdd FILL
XFILL_85_DFFSR_258 gnd vdd FILL
XFILL_20_DFFSR_180 gnd vdd FILL
XFILL_85_DFFSR_269 gnd vdd FILL
XFILL_20_DFFSR_191 gnd vdd FILL
XFILL_1_INVX1_120 gnd vdd FILL
XFILL_1_INVX1_131 gnd vdd FILL
XFILL_1_INVX1_142 gnd vdd FILL
XFILL_1_INVX1_153 gnd vdd FILL
XFILL_1_INVX1_164 gnd vdd FILL
XFILL_47_2_2 gnd vdd FILL
XFILL_1_INVX1_175 gnd vdd FILL
XFILL_8_NAND3X1_105 gnd vdd FILL
XFILL_8_NAND3X1_116 gnd vdd FILL
XFILL_1_INVX1_186 gnd vdd FILL
XFILL_1_INVX1_197 gnd vdd FILL
XFILL_24_DFFSR_190 gnd vdd FILL
XFILL_8_NAND3X1_127 gnd vdd FILL
XFILL_5_INVX1_130 gnd vdd FILL
XFILL_5_INVX1_141 gnd vdd FILL
XFILL_5_INVX1_152 gnd vdd FILL
XFILL_16_6_0 gnd vdd FILL
XFILL_5_INVX1_163 gnd vdd FILL
XFILL_5_INVX1_174 gnd vdd FILL
XFILL_5_INVX1_185 gnd vdd FILL
XFILL_5_INVX1_196 gnd vdd FILL
XFILL_30_1_2 gnd vdd FILL
XFILL_3_OAI22X1_3 gnd vdd FILL
XFILL_28_DFFSR_2 gnd vdd FILL
XFILL_85_DFFSR_3 gnd vdd FILL
XFILL_7_OAI22X1_2 gnd vdd FILL
XFILL_3_NAND3X1_101 gnd vdd FILL
XFILL_13_MUX2X1_140 gnd vdd FILL
XFILL_3_NAND3X1_112 gnd vdd FILL
XFILL_13_MUX2X1_151 gnd vdd FILL
XFILL_13_MUX2X1_162 gnd vdd FILL
XFILL_3_NAND3X1_123 gnd vdd FILL
XFILL_13_MUX2X1_173 gnd vdd FILL
XFILL_13_MUX2X1_184 gnd vdd FILL
XFILL_52_DFFSR_203 gnd vdd FILL
XFILL_52_DFFSR_214 gnd vdd FILL
XFILL_52_DFFSR_225 gnd vdd FILL
XFILL_52_DFFSR_236 gnd vdd FILL
XFILL_52_DFFSR_247 gnd vdd FILL
XFILL_52_DFFSR_258 gnd vdd FILL
XFILL_52_DFFSR_269 gnd vdd FILL
XFILL_66_5_0 gnd vdd FILL
XFILL_12_DFFSR_8 gnd vdd FILL
XFILL_38_2_2 gnd vdd FILL
XFILL_56_DFFSR_202 gnd vdd FILL
XFILL_29_CLKBUF1_19 gnd vdd FILL
XFILL_56_DFFSR_213 gnd vdd FILL
XFILL_56_DFFSR_224 gnd vdd FILL
XFILL_56_DFFSR_235 gnd vdd FILL
XFILL_56_DFFSR_246 gnd vdd FILL
XFILL_56_DFFSR_257 gnd vdd FILL
XFILL_56_DFFSR_268 gnd vdd FILL
XFILL_11_CLKBUF1_9 gnd vdd FILL
XFILL_83_DFFSR_102 gnd vdd FILL
XFILL_54_DFFSR_19 gnd vdd FILL
XFILL_83_DFFSR_113 gnd vdd FILL
XFILL_83_DFFSR_124 gnd vdd FILL
XFILL_83_DFFSR_135 gnd vdd FILL
XFILL_83_DFFSR_146 gnd vdd FILL
XFILL_83_DFFSR_157 gnd vdd FILL
XFILL_83_DFFSR_168 gnd vdd FILL
XFILL_83_DFFSR_179 gnd vdd FILL
XFILL_15_CLKBUF1_8 gnd vdd FILL
XFILL_3_DFFSR_205 gnd vdd FILL
XFILL_87_DFFSR_101 gnd vdd FILL
XFILL_3_DFFSR_216 gnd vdd FILL
XFILL_0_NAND3X1_5 gnd vdd FILL
XFILL_21_1_2 gnd vdd FILL
XFILL_87_DFFSR_112 gnd vdd FILL
XFILL_3_DFFSR_227 gnd vdd FILL
XFILL_87_DFFSR_123 gnd vdd FILL
XFILL_87_DFFSR_134 gnd vdd FILL
XFILL_3_DFFSR_238 gnd vdd FILL
XFILL_87_DFFSR_145 gnd vdd FILL
XFILL_3_DFFSR_249 gnd vdd FILL
XFILL_87_DFFSR_156 gnd vdd FILL
XFILL_11_BUFX4_103 gnd vdd FILL
XFILL_87_DFFSR_167 gnd vdd FILL
XFILL_14_BUFX4_50 gnd vdd FILL
XFILL_23_DFFSR_18 gnd vdd FILL
XFILL_23_DFFSR_29 gnd vdd FILL
XFILL_19_CLKBUF1_7 gnd vdd FILL
XFILL_87_DFFSR_178 gnd vdd FILL
XFILL_3_MUX2X1_190 gnd vdd FILL
XFILL_14_BUFX4_61 gnd vdd FILL
XFILL_87_DFFSR_189 gnd vdd FILL
XFILL_14_BUFX4_72 gnd vdd FILL
XFILL_7_DFFSR_204 gnd vdd FILL
XFILL_14_BUFX4_83 gnd vdd FILL
XFILL_7_DFFSR_215 gnd vdd FILL
XFILL_4_NAND3X1_4 gnd vdd FILL
XFILL_7_DFFSR_226 gnd vdd FILL
XDFFSR_240 INVX1_54/A DFFSR_52/CLK DFFSR_42/R vdd MUX2X1_41/Y gnd vdd DFFSR
XFILL_14_BUFX4_94 gnd vdd FILL
XFILL_7_DFFSR_237 gnd vdd FILL
XDFFSR_251 INVX1_48/A DFFSR_2/CLK BUFX4_50/Y vdd MUX2X1_34/Y gnd vdd DFFSR
XFILL_7_DFFSR_248 gnd vdd FILL
XDFFSR_262 NOR2X1_11/A DFFSR_1/CLK DFFSR_1/R vdd DFFSR_262/D gnd vdd DFFSR
XFILL_15_BUFX4_102 gnd vdd FILL
XFILL_63_DFFSR_17 gnd vdd FILL
XDFFSR_273 NOR2X1_5/A DFFSR_47/CLK DFFSR_26/R vdd DFFSR_273/D gnd vdd DFFSR
XFILL_7_DFFSR_259 gnd vdd FILL
XFILL_63_DFFSR_28 gnd vdd FILL
XFILL_63_DFFSR_39 gnd vdd FILL
XFILL_8_NAND3X1_3 gnd vdd FILL
XFILL_6_DFFSR_19 gnd vdd FILL
XFILL_32_DFFSR_16 gnd vdd FILL
XFILL_32_DFFSR_27 gnd vdd FILL
XFILL_32_DFFSR_38 gnd vdd FILL
XFILL_32_DFFSR_49 gnd vdd FILL
XFILL_57_5_0 gnd vdd FILL
XFILL_7_OAI22X1_17 gnd vdd FILL
XFILL_7_OAI22X1_28 gnd vdd FILL
XFILL_29_2_2 gnd vdd FILL
XFILL_4_2_2 gnd vdd FILL
XFILL_7_OAI22X1_39 gnd vdd FILL
XFILL_0_INVX1_209 gnd vdd FILL
XFILL_72_DFFSR_15 gnd vdd FILL
XFILL_23_DFFSR_202 gnd vdd FILL
XFILL_72_DFFSR_26 gnd vdd FILL
XFILL_23_DFFSR_213 gnd vdd FILL
XFILL_72_DFFSR_37 gnd vdd FILL
XFILL_23_DFFSR_224 gnd vdd FILL
XFILL_15_MUX2X1_5 gnd vdd FILL
XFILL_72_DFFSR_48 gnd vdd FILL
XFILL_4_AOI22X1_9 gnd vdd FILL
XFILL_23_DFFSR_235 gnd vdd FILL
XFILL_72_DFFSR_59 gnd vdd FILL
XFILL_23_DFFSR_246 gnd vdd FILL
XFILL_23_DFFSR_257 gnd vdd FILL
XFILL_23_DFFSR_268 gnd vdd FILL
XFILL_6_NAND3X1_60 gnd vdd FILL
XFILL_6_NAND3X1_71 gnd vdd FILL
XFILL_4_INVX1_208 gnd vdd FILL
XFILL_50_DFFSR_102 gnd vdd FILL
XFILL_6_NAND3X1_82 gnd vdd FILL
XFILL_27_DFFSR_201 gnd vdd FILL
XFILL_6_NAND3X1_93 gnd vdd FILL
XFILL_4_INVX1_219 gnd vdd FILL
XFILL_27_DFFSR_212 gnd vdd FILL
XFILL_50_DFFSR_113 gnd vdd FILL
XFILL_50_DFFSR_124 gnd vdd FILL
XFILL_27_DFFSR_223 gnd vdd FILL
XFILL_27_DFFSR_234 gnd vdd FILL
XFILL_6_BUFX4_60 gnd vdd FILL
XFILL_50_DFFSR_135 gnd vdd FILL
XFILL_8_AOI22X1_8 gnd vdd FILL
XFILL_50_DFFSR_146 gnd vdd FILL
XFILL_40_4_0 gnd vdd FILL
XFILL_41_DFFSR_14 gnd vdd FILL
XFILL_6_BUFX4_71 gnd vdd FILL
XFILL_41_DFFSR_25 gnd vdd FILL
XFILL_27_DFFSR_245 gnd vdd FILL
XFILL_12_1_2 gnd vdd FILL
XFILL_50_DFFSR_157 gnd vdd FILL
XFILL_41_DFFSR_36 gnd vdd FILL
XFILL_27_DFFSR_256 gnd vdd FILL
XFILL_6_BUFX4_82 gnd vdd FILL
XFILL_6_BUFX4_93 gnd vdd FILL
XFILL_27_DFFSR_267 gnd vdd FILL
XFILL_50_DFFSR_168 gnd vdd FILL
XFILL_41_DFFSR_47 gnd vdd FILL
XFILL_50_DFFSR_179 gnd vdd FILL
XFILL_54_DFFSR_101 gnd vdd FILL
XFILL_41_DFFSR_58 gnd vdd FILL
XFILL_0_OAI21X1_19 gnd vdd FILL
XFILL_8_BUFX2_1 gnd vdd FILL
XFILL_41_DFFSR_69 gnd vdd FILL
XFILL_18_CLKBUF1_15 gnd vdd FILL
XFILL_54_DFFSR_112 gnd vdd FILL
XFILL_18_CLKBUF1_26 gnd vdd FILL
XFILL_54_DFFSR_123 gnd vdd FILL
XFILL_54_DFFSR_134 gnd vdd FILL
XFILL_18_CLKBUF1_37 gnd vdd FILL
XFILL_81_DFFSR_13 gnd vdd FILL
XFILL_54_DFFSR_145 gnd vdd FILL
XFILL_13_AOI21X1_12 gnd vdd FILL
XFILL_54_DFFSR_156 gnd vdd FILL
XFILL_81_DFFSR_24 gnd vdd FILL
XFILL_81_DFFSR_35 gnd vdd FILL
XFILL_13_AOI21X1_23 gnd vdd FILL
XFILL_13_AOI21X1_34 gnd vdd FILL
XFILL_81_DFFSR_46 gnd vdd FILL
XFILL_54_DFFSR_167 gnd vdd FILL
XFILL_13_AOI21X1_45 gnd vdd FILL
XFILL_54_DFFSR_178 gnd vdd FILL
XFILL_81_DFFSR_57 gnd vdd FILL
XFILL_10_DFFSR_13 gnd vdd FILL
XFILL_58_DFFSR_100 gnd vdd FILL
XFILL_54_DFFSR_189 gnd vdd FILL
XFILL_13_AOI21X1_56 gnd vdd FILL
XFILL_81_DFFSR_68 gnd vdd FILL
XFILL_10_DFFSR_24 gnd vdd FILL
XFILL_58_DFFSR_111 gnd vdd FILL
XFILL_13_AOI21X1_67 gnd vdd FILL
XFILL_10_DFFSR_35 gnd vdd FILL
XFILL_81_DFFSR_79 gnd vdd FILL
XFILL_13_AOI21X1_78 gnd vdd FILL
XFILL_10_DFFSR_46 gnd vdd FILL
XFILL_58_DFFSR_122 gnd vdd FILL
XFILL_58_DFFSR_133 gnd vdd FILL
XFILL_10_DFFSR_57 gnd vdd FILL
XFILL_58_DFFSR_144 gnd vdd FILL
XFILL_8_NOR2X1_6 gnd vdd FILL
XFILL_58_DFFSR_155 gnd vdd FILL
XFILL_10_DFFSR_68 gnd vdd FILL
XFILL_10_DFFSR_79 gnd vdd FILL
XFILL_58_DFFSR_166 gnd vdd FILL
XFILL_1_DFFSR_104 gnd vdd FILL
XFILL_58_DFFSR_177 gnd vdd FILL
XFILL_50_DFFSR_12 gnd vdd FILL
XFILL_58_DFFSR_188 gnd vdd FILL
XFILL_1_DFFSR_115 gnd vdd FILL
XFILL_58_DFFSR_199 gnd vdd FILL
XFILL_50_DFFSR_23 gnd vdd FILL
XFILL_1_DFFSR_126 gnd vdd FILL
XFILL_50_DFFSR_34 gnd vdd FILL
XFILL_1_DFFSR_137 gnd vdd FILL
XFILL_21_NOR3X1_9 gnd vdd FILL
XFILL_50_DFFSR_45 gnd vdd FILL
XFILL_50_DFFSR_56 gnd vdd FILL
XFILL_1_DFFSR_148 gnd vdd FILL
XFILL_50_DFFSR_67 gnd vdd FILL
XFILL_1_DFFSR_159 gnd vdd FILL
XFILL_50_DFFSR_78 gnd vdd FILL
XFILL_50_DFFSR_89 gnd vdd FILL
XFILL_5_DFFSR_103 gnd vdd FILL
XFILL_48_5_0 gnd vdd FILL
XFILL_5_DFFSR_114 gnd vdd FILL
XFILL_7_MUX2X1_4 gnd vdd FILL
XFILL_5_DFFSR_125 gnd vdd FILL
XFILL_5_DFFSR_136 gnd vdd FILL
XFILL_5_DFFSR_147 gnd vdd FILL
XFILL_5_DFFSR_158 gnd vdd FILL
XFILL_51_DFFSR_6 gnd vdd FILL
XFILL_5_DFFSR_169 gnd vdd FILL
XFILL_9_NAND3X1_106 gnd vdd FILL
XFILL_9_DFFSR_102 gnd vdd FILL
XFILL_9_NAND3X1_117 gnd vdd FILL
XFILL_8_CLKBUF1_10 gnd vdd FILL
XFILL_8_CLKBUF1_21 gnd vdd FILL
XFILL_13_MUX2X1_11 gnd vdd FILL
XFILL_9_DFFSR_113 gnd vdd FILL
XFILL_8_CLKBUF1_32 gnd vdd FILL
XFILL_9_NAND3X1_128 gnd vdd FILL
XFILL_9_DFFSR_124 gnd vdd FILL
XFILL_62_0_2 gnd vdd FILL
XFILL_13_MUX2X1_22 gnd vdd FILL
XFILL_9_DFFSR_135 gnd vdd FILL
XFILL_16_MUX2X1_106 gnd vdd FILL
XFILL_13_MUX2X1_33 gnd vdd FILL
XFILL_9_DFFSR_146 gnd vdd FILL
XFILL_13_MUX2X1_44 gnd vdd FILL
XFILL_9_DFFSR_157 gnd vdd FILL
XFILL_16_MUX2X1_117 gnd vdd FILL
XFILL_13_MUX2X1_55 gnd vdd FILL
XFILL_13_MUX2X1_66 gnd vdd FILL
XFILL_9_DFFSR_168 gnd vdd FILL
XFILL_16_MUX2X1_128 gnd vdd FILL
XFILL_3_AOI21X1_40 gnd vdd FILL
XFILL_16_MUX2X1_139 gnd vdd FILL
XFILL_30_NOR3X1_7 gnd vdd FILL
XFILL_13_MUX2X1_77 gnd vdd FILL
XFILL_9_DFFSR_179 gnd vdd FILL
XFILL_3_AOI21X1_51 gnd vdd FILL
XFILL_1_NOR3X1_15 gnd vdd FILL
XFILL_13_MUX2X1_88 gnd vdd FILL
XFILL_1_NOR3X1_26 gnd vdd FILL
XOAI21X1_10 INVX1_31/Y NOR2X1_51/B OAI21X1_10/C gnd NOR2X1_67/A vdd OAI21X1
XFILL_3_AOI21X1_62 gnd vdd FILL
XFILL_13_MUX2X1_99 gnd vdd FILL
XOAI21X1_21 INVX1_157/Y OAI21X1_3/B OAI21X1_21/C gnd NOR2X1_92/A vdd OAI21X1
XFILL_3_AOI21X1_73 gnd vdd FILL
XFILL_17_MUX2X1_10 gnd vdd FILL
XFILL_13_OAI22X1_20 gnd vdd FILL
XFILL_17_MUX2X1_21 gnd vdd FILL
XFILL_13_OAI22X1_31 gnd vdd FILL
XOAI21X1_32 INVX1_191/Y OAI21X1_7/B OAI21X1_32/C gnd OAI21X1_32/Y vdd OAI21X1
XFILL_31_4_0 gnd vdd FILL
XFILL_1_NOR3X1_37 gnd vdd FILL
XFILL_13_OAI22X1_42 gnd vdd FILL
XOAI21X1_43 OAI21X1_1/A OAI21X1_1/B INVX2_4/A gnd OAI21X1_43/Y vdd OAI21X1
XFILL_1_NOR3X1_48 gnd vdd FILL
XFILL_17_MUX2X1_32 gnd vdd FILL
XFILL_17_MUX2X1_43 gnd vdd FILL
XFILL_17_MUX2X1_54 gnd vdd FILL
XFILL_2_DFFSR_12 gnd vdd FILL
XFILL_17_MUX2X1_65 gnd vdd FILL
XFILL_2_DFFSR_23 gnd vdd FILL
XFILL_5_NOR3X1_14 gnd vdd FILL
XFILL_17_MUX2X1_76 gnd vdd FILL
XFILL_6_NOR2X1_150 gnd vdd FILL
XFILL_17_MUX2X1_87 gnd vdd FILL
XFILL_6_NOR2X1_161 gnd vdd FILL
XFILL_2_DFFSR_34 gnd vdd FILL
XFILL_5_NOR3X1_25 gnd vdd FILL
XFILL_16_DFFSR_9 gnd vdd FILL
XFILL_5_NOR3X1_36 gnd vdd FILL
XFILL_2_DFFSR_45 gnd vdd FILL
XFILL_13_NAND3X1_130 gnd vdd FILL
XFILL_17_MUX2X1_98 gnd vdd FILL
XFILL_6_NOR2X1_172 gnd vdd FILL
XFILL_2_DFFSR_56 gnd vdd FILL
XFILL_21_DFFSR_101 gnd vdd FILL
XFILL_5_NOR3X1_47 gnd vdd FILL
XFILL_2_DFFSR_67 gnd vdd FILL
XFILL_6_NOR2X1_183 gnd vdd FILL
XFILL_2_DFFSR_78 gnd vdd FILL
XFILL_6_NOR2X1_194 gnd vdd FILL
XFILL_21_DFFSR_112 gnd vdd FILL
XFILL_21_DFFSR_123 gnd vdd FILL
XFILL_2_DFFSR_89 gnd vdd FILL
XFILL_21_DFFSR_134 gnd vdd FILL
XFILL_21_DFFSR_145 gnd vdd FILL
XFILL_10_NOR2X1_200 gnd vdd FILL
XFILL_21_DFFSR_156 gnd vdd FILL
XFILL_9_NOR3X1_13 gnd vdd FILL
XFILL_9_NOR3X1_24 gnd vdd FILL
XFILL_21_DFFSR_167 gnd vdd FILL
XFILL_21_DFFSR_178 gnd vdd FILL
XFILL_2_INVX1_107 gnd vdd FILL
XFILL_9_NOR3X1_35 gnd vdd FILL
XFILL_9_NOR3X1_46 gnd vdd FILL
XFILL_25_DFFSR_100 gnd vdd FILL
XFILL_21_DFFSR_189 gnd vdd FILL
XFILL_2_INVX1_118 gnd vdd FILL
XFILL_25_DFFSR_111 gnd vdd FILL
XFILL_2_INVX1_129 gnd vdd FILL
XFILL_25_DFFSR_122 gnd vdd FILL
XFILL_25_DFFSR_133 gnd vdd FILL
XFILL_25_DFFSR_144 gnd vdd FILL
XFILL_25_DFFSR_155 gnd vdd FILL
XFILL_4_NAND3X1_102 gnd vdd FILL
XFILL_23_MUX2X1_130 gnd vdd FILL
XFILL_4_NAND3X1_113 gnd vdd FILL
XFILL_23_MUX2X1_141 gnd vdd FILL
XFILL_25_DFFSR_166 gnd vdd FILL
XFILL_23_MUX2X1_152 gnd vdd FILL
XFILL_23_MUX2X1_163 gnd vdd FILL
XFILL_25_DFFSR_177 gnd vdd FILL
XFILL_6_INVX1_106 gnd vdd FILL
XFILL_4_NAND3X1_124 gnd vdd FILL
XFILL_25_DFFSR_188 gnd vdd FILL
XFILL_6_MUX2X1_101 gnd vdd FILL
XFILL_6_INVX1_117 gnd vdd FILL
XFILL_6_MUX2X1_112 gnd vdd FILL
XFILL_29_DFFSR_110 gnd vdd FILL
XFILL_25_DFFSR_199 gnd vdd FILL
XFILL_23_MUX2X1_174 gnd vdd FILL
XFILL_6_MUX2X1_123 gnd vdd FILL
XFILL_23_MUX2X1_185 gnd vdd FILL
XFILL_6_INVX1_128 gnd vdd FILL
XFILL_29_DFFSR_121 gnd vdd FILL
XFILL_6_INVX1_139 gnd vdd FILL
XFILL_6_MUX2X1_134 gnd vdd FILL
XFILL_29_DFFSR_132 gnd vdd FILL
XFILL_6_MUX2X1_145 gnd vdd FILL
XFILL_29_DFFSR_143 gnd vdd FILL
XFILL_29_DFFSR_154 gnd vdd FILL
XFILL_6_MUX2X1_156 gnd vdd FILL
XFILL_39_5_0 gnd vdd FILL
XFILL_29_DFFSR_165 gnd vdd FILL
XFILL_6_MUX2X1_167 gnd vdd FILL
XFILL_6_MUX2X1_178 gnd vdd FILL
XFILL_21_NOR3X1_12 gnd vdd FILL
XFILL_29_DFFSR_176 gnd vdd FILL
XFILL_19_DFFSR_90 gnd vdd FILL
XFILL_6_MUX2X1_189 gnd vdd FILL
XFILL_29_DFFSR_187 gnd vdd FILL
XFILL_21_NOR3X1_23 gnd vdd FILL
XFILL_21_NOR3X1_34 gnd vdd FILL
XFILL_29_DFFSR_198 gnd vdd FILL
XFILL_71_DFFSR_201 gnd vdd FILL
XFILL_21_NOR3X1_45 gnd vdd FILL
XFILL_71_DFFSR_212 gnd vdd FILL
XFILL_7_OAI21X1_50 gnd vdd FILL
XFILL_71_DFFSR_223 gnd vdd FILL
XFILL_71_DFFSR_234 gnd vdd FILL
XFILL_53_0_2 gnd vdd FILL
XFILL_71_DFFSR_245 gnd vdd FILL
XFILL_25_NOR3X1_11 gnd vdd FILL
XFILL_71_DFFSR_256 gnd vdd FILL
XFILL_71_DFFSR_267 gnd vdd FILL
XFILL_25_NOR3X1_22 gnd vdd FILL
XFILL_25_NOR3X1_33 gnd vdd FILL
XFILL_25_NOR3X1_44 gnd vdd FILL
XFILL_75_DFFSR_200 gnd vdd FILL
XFILL_75_DFFSR_211 gnd vdd FILL
XFILL_75_DFFSR_222 gnd vdd FILL
XFILL_75_DFFSR_233 gnd vdd FILL
XFILL_22_4_0 gnd vdd FILL
XFILL_10_BUFX4_9 gnd vdd FILL
XFILL_75_DFFSR_244 gnd vdd FILL
XFILL_29_NOR3X1_10 gnd vdd FILL
XFILL_75_DFFSR_255 gnd vdd FILL
XFILL_75_DFFSR_266 gnd vdd FILL
XFILL_29_NOR3X1_21 gnd vdd FILL
XFILL_30_CLKBUF1_7 gnd vdd FILL
XFILL_29_NOR3X1_32 gnd vdd FILL
XFILL_29_NOR3X1_43 gnd vdd FILL
XFILL_79_DFFSR_210 gnd vdd FILL
XFILL_79_DFFSR_221 gnd vdd FILL
XFILL_79_DFFSR_232 gnd vdd FILL
XFILL_79_DFFSR_243 gnd vdd FILL
XFILL_79_DFFSR_254 gnd vdd FILL
XFILL_79_DFFSR_265 gnd vdd FILL
XFILL_34_CLKBUF1_6 gnd vdd FILL
XFILL_9_NAND3X1_15 gnd vdd FILL
XFILL_9_NAND3X1_26 gnd vdd FILL
XFILL_9_NAND3X1_37 gnd vdd FILL
XFILL_9_NAND3X1_48 gnd vdd FILL
XFILL_9_NAND3X1_59 gnd vdd FILL
XFILL_15_BUFX4_17 gnd vdd FILL
XFILL_15_BUFX4_28 gnd vdd FILL
XFILL_0_NOR3X1_3 gnd vdd FILL
XFILL_15_BUFX4_39 gnd vdd FILL
XFILL_5_5_0 gnd vdd FILL
XFILL_2_NAND2X1_17 gnd vdd FILL
XFILL_33_DFFSR_3 gnd vdd FILL
XFILL_2_NAND2X1_28 gnd vdd FILL
XFILL_2_NAND2X1_39 gnd vdd FILL
XFILL_44_0_2 gnd vdd FILL
XFILL_0_OAI21X1_2 gnd vdd FILL
XFILL_12_MUX2X1_170 gnd vdd FILL
XFILL_13_4_0 gnd vdd FILL
XFILL_12_MUX2X1_181 gnd vdd FILL
XFILL_42_DFFSR_200 gnd vdd FILL
XFILL_12_MUX2X1_192 gnd vdd FILL
XFILL_42_DFFSR_211 gnd vdd FILL
XFILL_42_DFFSR_222 gnd vdd FILL
XFILL_4_OAI21X1_1 gnd vdd FILL
XFILL_42_DFFSR_233 gnd vdd FILL
XFILL_42_DFFSR_244 gnd vdd FILL
XFILL_42_DFFSR_255 gnd vdd FILL
XFILL_1_NOR2X1_70 gnd vdd FILL
XFILL_42_DFFSR_266 gnd vdd FILL
XFILL_1_NOR2X1_81 gnd vdd FILL
XFILL_1_NOR2X1_92 gnd vdd FILL
XFILL_28_CLKBUF1_16 gnd vdd FILL
XFILL_46_DFFSR_210 gnd vdd FILL
XFILL_46_DFFSR_221 gnd vdd FILL
XFILL_28_CLKBUF1_27 gnd vdd FILL
XFILL_28_CLKBUF1_38 gnd vdd FILL
XFILL_46_DFFSR_232 gnd vdd FILL
XFILL_55_DFFSR_7 gnd vdd FILL
XFILL_7_BUFX4_16 gnd vdd FILL
XFILL_46_DFFSR_243 gnd vdd FILL
XFILL_7_BUFX4_27 gnd vdd FILL
XFILL_46_DFFSR_254 gnd vdd FILL
XFILL_7_BUFX4_38 gnd vdd FILL
XFILL_5_NOR2X1_80 gnd vdd FILL
XFILL_7_BUFX4_49 gnd vdd FILL
XFILL_46_DFFSR_265 gnd vdd FILL
XFILL_5_NOR2X1_91 gnd vdd FILL
XFILL_73_DFFSR_110 gnd vdd FILL
XFILL_6_AOI21X1_17 gnd vdd FILL
XFILL_73_DFFSR_121 gnd vdd FILL
XFILL_73_DFFSR_132 gnd vdd FILL
XFILL_6_AOI21X1_28 gnd vdd FILL
XFILL_73_DFFSR_143 gnd vdd FILL
XFILL_73_DFFSR_154 gnd vdd FILL
XFILL_6_AOI21X1_39 gnd vdd FILL
XFILL_73_DFFSR_165 gnd vdd FILL
XFILL_16_OAI22X1_19 gnd vdd FILL
XFILL_73_DFFSR_176 gnd vdd FILL
XFILL_9_NOR2X1_90 gnd vdd FILL
XFILL_73_DFFSR_187 gnd vdd FILL
XFILL_6_3 gnd vdd FILL
XFILL_73_DFFSR_198 gnd vdd FILL
XFILL_9_NOR2X1_105 gnd vdd FILL
XFILL_77_DFFSR_120 gnd vdd FILL
XFILL_9_NOR2X1_116 gnd vdd FILL
XFILL_77_DFFSR_131 gnd vdd FILL
XFILL_77_DFFSR_142 gnd vdd FILL
XFILL_9_NOR2X1_127 gnd vdd FILL
XFILL_62_5 gnd vdd FILL
XFILL_77_DFFSR_153 gnd vdd FILL
XFILL_9_NOR2X1_138 gnd vdd FILL
XFILL_9_NOR2X1_149 gnd vdd FILL
XFILL_77_DFFSR_164 gnd vdd FILL
XFILL_77_DFFSR_175 gnd vdd FILL
XFILL_15_NAND3X1_40 gnd vdd FILL
XFILL_77_DFFSR_186 gnd vdd FILL
XFILL_15_NAND3X1_51 gnd vdd FILL
XFILL_15_NAND3X1_62 gnd vdd FILL
XFILL_77_DFFSR_197 gnd vdd FILL
XFILL_14_AND2X2_4 gnd vdd FILL
XFILL_15_NAND3X1_73 gnd vdd FILL
XFILL_15_NAND3X1_84 gnd vdd FILL
XFILL_15_NAND3X1_95 gnd vdd FILL
XFILL_35_CLKBUF1_40 gnd vdd FILL
XFILL_63_3_0 gnd vdd FILL
XFILL_35_0_2 gnd vdd FILL
XFILL_1_NAND2X1_3 gnd vdd FILL
XFILL_11_BUFX4_10 gnd vdd FILL
XFILL_11_BUFX4_21 gnd vdd FILL
XFILL_11_BUFX4_32 gnd vdd FILL
XFILL_11_BUFX4_43 gnd vdd FILL
XFILL_5_NAND2X1_2 gnd vdd FILL
XFILL_59_DFFSR_109 gnd vdd FILL
XFILL_11_BUFX4_54 gnd vdd FILL
XFILL_11_BUFX4_65 gnd vdd FILL
XFILL_11_BUFX4_76 gnd vdd FILL
XFILL_11_BUFX4_87 gnd vdd FILL
XFILL_6_OAI22X1_14 gnd vdd FILL
XFILL_11_BUFX4_98 gnd vdd FILL
XFILL_6_OAI22X1_25 gnd vdd FILL
XFILL_6_OAI22X1_36 gnd vdd FILL
XDFFSR_13 DFFSR_13/Q DFFSR_97/CLK DFFSR_97/R vdd DFFSR_13/D gnd vdd DFFSR
XFILL_14_NAND3X1_120 gnd vdd FILL
XFILL_14_NAND3X1_131 gnd vdd FILL
XFILL_6_OAI22X1_47 gnd vdd FILL
XFILL_9_NAND2X1_1 gnd vdd FILL
XDFFSR_24 DFFSR_24/Q CLKBUF1_8/Y DFFSR_55/R vdd DFFSR_24/D gnd vdd DFFSR
XDFFSR_35 DFFSR_35/Q DFFSR_81/CLK DFFSR_53/R vdd DFFSR_35/D gnd vdd DFFSR
XFILL_13_DFFSR_210 gnd vdd FILL
XDFFSR_46 DFFSR_46/Q DFFSR_78/CLK DFFSR_78/R vdd DFFSR_46/D gnd vdd DFFSR
XDFFSR_57 DFFSR_57/Q DFFSR_57/CLK DFFSR_57/R vdd DFFSR_57/D gnd vdd DFFSR
XFILL_13_DFFSR_221 gnd vdd FILL
XFILL_13_DFFSR_232 gnd vdd FILL
XDFFSR_68 DFFSR_68/Q DFFSR_90/CLK DFFSR_90/R vdd DFFSR_68/D gnd vdd DFFSR
XFILL_13_DFFSR_243 gnd vdd FILL
XDFFSR_79 DFFSR_79/Q DFFSR_79/CLK DFFSR_79/R vdd DFFSR_79/D gnd vdd DFFSR
XFILL_13_DFFSR_254 gnd vdd FILL
XFILL_13_DFFSR_265 gnd vdd FILL
XFILL_40_DFFSR_110 gnd vdd FILL
XFILL_5_NAND3X1_90 gnd vdd FILL
XFILL_3_NOR2X1_205 gnd vdd FILL
XFILL_17_DFFSR_220 gnd vdd FILL
XFILL_40_DFFSR_121 gnd vdd FILL
XFILL_40_DFFSR_132 gnd vdd FILL
XFILL_1_AOI21X1_8 gnd vdd FILL
XFILL_9_NAND2X1_70 gnd vdd FILL
XFILL_17_DFFSR_231 gnd vdd FILL
XFILL_5_INVX1_11 gnd vdd FILL
XFILL_40_DFFSR_143 gnd vdd FILL
XFILL_9_NAND2X1_81 gnd vdd FILL
XFILL_5_INVX1_22 gnd vdd FILL
XFILL_40_DFFSR_154 gnd vdd FILL
XCLKBUF1_11 BUFX4_84/Y gnd DFFSR_70/CLK vdd CLKBUF1
XFILL_17_DFFSR_242 gnd vdd FILL
XFILL_5_NAND3X1_103 gnd vdd FILL
XFILL_9_NAND2X1_92 gnd vdd FILL
XCLKBUF1_22 BUFX4_4/Y gnd DFFSR_8/CLK vdd CLKBUF1
XFILL_5_NAND3X1_114 gnd vdd FILL
XFILL_17_DFFSR_253 gnd vdd FILL
XFILL_5_INVX1_33 gnd vdd FILL
XFILL_40_DFFSR_165 gnd vdd FILL
XCLKBUF1_33 BUFX4_95/Y gnd DFFSR_79/CLK vdd CLKBUF1
XFILL_5_NAND3X1_125 gnd vdd FILL
XFILL_5_INVX1_44 gnd vdd FILL
XFILL_17_DFFSR_264 gnd vdd FILL
XFILL_6_AND2X2_3 gnd vdd FILL
XFILL_17_DFFSR_275 gnd vdd FILL
XFILL_5_INVX1_55 gnd vdd FILL
XFILL_40_DFFSR_176 gnd vdd FILL
XFILL_5_INVX1_66 gnd vdd FILL
XFILL_40_DFFSR_187 gnd vdd FILL
XFILL_17_CLKBUF1_12 gnd vdd FILL
XFILL_5_INVX1_77 gnd vdd FILL
XFILL_40_DFFSR_198 gnd vdd FILL
XFILL_17_CLKBUF1_23 gnd vdd FILL
XFILL_5_INVX1_88 gnd vdd FILL
XFILL_44_DFFSR_120 gnd vdd FILL
XFILL_44_DFFSR_131 gnd vdd FILL
XFILL_5_AOI21X1_7 gnd vdd FILL
XFILL_17_CLKBUF1_34 gnd vdd FILL
XFILL_5_INVX1_99 gnd vdd FILL
XFILL_44_DFFSR_142 gnd vdd FILL
XFILL_44_DFFSR_153 gnd vdd FILL
XFILL_12_AOI21X1_20 gnd vdd FILL
XFILL_44_DFFSR_164 gnd vdd FILL
XFILL_12_AOI21X1_31 gnd vdd FILL
XFILL_12_MUX2X1_9 gnd vdd FILL
XFILL_12_AOI21X1_42 gnd vdd FILL
XFILL_44_DFFSR_175 gnd vdd FILL
XFILL_2_DFFSR_2 gnd vdd FILL
XFILL_18_MUX2X1_19 gnd vdd FILL
XFILL_44_DFFSR_186 gnd vdd FILL
XFILL_12_AOI21X1_53 gnd vdd FILL
XFILL_54_3_0 gnd vdd FILL
XFILL_44_DFFSR_197 gnd vdd FILL
XFILL_12_AOI21X1_64 gnd vdd FILL
XFILL_1_0_2 gnd vdd FILL
XFILL_12_AOI21X1_75 gnd vdd FILL
XFILL_26_0_2 gnd vdd FILL
XFILL_48_DFFSR_130 gnd vdd FILL
XFILL_3_BUFX4_20 gnd vdd FILL
XFILL_9_AOI21X1_6 gnd vdd FILL
XFILL_72_DFFSR_1 gnd vdd FILL
XFILL_3_BUFX4_31 gnd vdd FILL
XFILL_48_DFFSR_141 gnd vdd FILL
XFILL_48_DFFSR_152 gnd vdd FILL
XFILL_3_BUFX4_42 gnd vdd FILL
XFILL_10_AOI22X1_4 gnd vdd FILL
XFILL_3_BUFX4_53 gnd vdd FILL
XFILL_48_DFFSR_163 gnd vdd FILL
XFILL_48_DFFSR_174 gnd vdd FILL
XFILL_3_BUFX4_64 gnd vdd FILL
XFILL_48_DFFSR_185 gnd vdd FILL
XFILL_3_BUFX4_75 gnd vdd FILL
XFILL_3_BUFX4_86 gnd vdd FILL
XFILL_48_DFFSR_196 gnd vdd FILL
XFILL_3_BUFX4_97 gnd vdd FILL
XFILL_10_BUFX2_6 gnd vdd FILL
XFILL_14_AOI22X1_3 gnd vdd FILL
XFILL_26_DFFSR_109 gnd vdd FILL
XFILL_21_MUX2X1_7 gnd vdd FILL
XFILL_18_AOI22X1_2 gnd vdd FILL
XFILL_0_NAND3X1_110 gnd vdd FILL
XFILL_0_NAND3X1_121 gnd vdd FILL
XFILL_37_DFFSR_4 gnd vdd FILL
XINVX1_107 INVX1_107/A gnd MUX2X1_94/A vdd INVX1
XINVX1_118 DFFSR_46/Q gnd NOR3X1_46/A vdd INVX1
XFILL_0_NAND3X1_132 gnd vdd FILL
XINVX1_129 INVX1_129/A gnd INVX1_129/Y vdd INVX1
XFILL_29_DFFSR_11 gnd vdd FILL
XFILL_29_DFFSR_22 gnd vdd FILL
XFILL_7_CLKBUF1_40 gnd vdd FILL
XFILL_15_MUX2X1_103 gnd vdd FILL
XFILL_15_MUX2X1_114 gnd vdd FILL
XFILL_29_DFFSR_33 gnd vdd FILL
XFILL_29_DFFSR_44 gnd vdd FILL
XFILL_15_MUX2X1_125 gnd vdd FILL
XFILL_29_DFFSR_55 gnd vdd FILL
XFILL_29_DFFSR_66 gnd vdd FILL
XFILL_15_MUX2X1_136 gnd vdd FILL
XFILL_29_DFFSR_77 gnd vdd FILL
XFILL_15_MUX2X1_147 gnd vdd FILL
XFILL_15_MUX2X1_158 gnd vdd FILL
XFILL_9_1_2 gnd vdd FILL
XFILL_2_AOI21X1_70 gnd vdd FILL
XFILL_15_MUX2X1_169 gnd vdd FILL
XFILL_29_DFFSR_88 gnd vdd FILL
XFILL_2_AOI21X1_81 gnd vdd FILL
XFILL_29_DFFSR_99 gnd vdd FILL
XFILL_69_DFFSR_10 gnd vdd FILL
XFILL_69_DFFSR_21 gnd vdd FILL
XFILL_12_OAI22X1_50 gnd vdd FILL
XFILL_69_DFFSR_32 gnd vdd FILL
XFILL_69_DFFSR_43 gnd vdd FILL
XFILL_4_MUX2X1_8 gnd vdd FILL
XFILL_69_DFFSR_54 gnd vdd FILL
XFILL_69_DFFSR_65 gnd vdd FILL
XFILL_69_DFFSR_76 gnd vdd FILL
XFILL_69_DFFSR_87 gnd vdd FILL
XFILL_69_DFFSR_98 gnd vdd FILL
XFILL_5_NOR2X1_180 gnd vdd FILL
XFILL_5_NOR2X1_191 gnd vdd FILL
XFILL_11_DFFSR_120 gnd vdd FILL
XFILL_76_DFFSR_209 gnd vdd FILL
XFILL_11_DFFSR_131 gnd vdd FILL
XFILL_59_DFFSR_8 gnd vdd FILL
XFILL_11_DFFSR_142 gnd vdd FILL
XFILL_11_DFFSR_153 gnd vdd FILL
XFILL_38_DFFSR_20 gnd vdd FILL
XFILL_45_3_0 gnd vdd FILL
XFILL_38_DFFSR_31 gnd vdd FILL
XFILL_11_DFFSR_164 gnd vdd FILL
XFILL_38_DFFSR_42 gnd vdd FILL
XFILL_17_0_2 gnd vdd FILL
XFILL_0_CLKBUF1_7 gnd vdd FILL
XFILL_11_DFFSR_175 gnd vdd FILL
XFILL_11_DFFSR_186 gnd vdd FILL
XFILL_38_DFFSR_53 gnd vdd FILL
XFILL_11_DFFSR_197 gnd vdd FILL
XFILL_38_DFFSR_64 gnd vdd FILL
XFILL_38_DFFSR_75 gnd vdd FILL
XFILL_38_DFFSR_86 gnd vdd FILL
XFILL_15_DFFSR_130 gnd vdd FILL
XFILL_38_DFFSR_97 gnd vdd FILL
XFILL_15_DFFSR_141 gnd vdd FILL
XFILL_15_DFFSR_152 gnd vdd FILL
XFILL_27_8 gnd vdd FILL
XFILL_78_DFFSR_30 gnd vdd FILL
XFILL_15_DFFSR_163 gnd vdd FILL
XFILL_78_DFFSR_41 gnd vdd FILL
XFILL_15_DFFSR_174 gnd vdd FILL
XFILL_22_MUX2X1_160 gnd vdd FILL
XFILL_78_DFFSR_52 gnd vdd FILL
XFILL_4_CLKBUF1_6 gnd vdd FILL
XFILL_22_MUX2X1_171 gnd vdd FILL
XFILL_15_DFFSR_185 gnd vdd FILL
XFILL_78_DFFSR_63 gnd vdd FILL
XFILL_15_DFFSR_196 gnd vdd FILL
XFILL_5_MUX2X1_120 gnd vdd FILL
XFILL_78_DFFSR_74 gnd vdd FILL
XFILL_22_MUX2X1_182 gnd vdd FILL
XFILL_78_DFFSR_85 gnd vdd FILL
XFILL_5_MUX2X1_131 gnd vdd FILL
XFILL_22_MUX2X1_193 gnd vdd FILL
XFILL_78_DFFSR_96 gnd vdd FILL
XFILL_5_MUX2X1_142 gnd vdd FILL
XFILL_19_DFFSR_140 gnd vdd FILL
XFILL_5_MUX2X1_153 gnd vdd FILL
XFILL_0_BUFX4_101 gnd vdd FILL
XFILL_19_DFFSR_151 gnd vdd FILL
XFILL_19_DFFSR_162 gnd vdd FILL
XFILL_5_MUX2X1_164 gnd vdd FILL
XFILL_5_MUX2X1_175 gnd vdd FILL
XFILL_19_DFFSR_173 gnd vdd FILL
XFILL_5_MUX2X1_186 gnd vdd FILL
XFILL_1_INVX1_70 gnd vdd FILL
XFILL_8_CLKBUF1_5 gnd vdd FILL
XFILL_19_DFFSR_184 gnd vdd FILL
XFILL_1_INVX1_81 gnd vdd FILL
XFILL_11_NOR3X1_20 gnd vdd FILL
XFILL_1_INVX1_92 gnd vdd FILL
XFILL_11_NOR3X1_31 gnd vdd FILL
XFILL_19_DFFSR_195 gnd vdd FILL
XFILL_11_NOR3X1_42 gnd vdd FILL
XFILL_47_DFFSR_40 gnd vdd FILL
XFILL_18_NOR3X1_4 gnd vdd FILL
XFILL_47_DFFSR_51 gnd vdd FILL
XFILL_47_DFFSR_62 gnd vdd FILL
XFILL_61_DFFSR_220 gnd vdd FILL
XFILL_61_DFFSR_231 gnd vdd FILL
XFILL_4_BUFX4_100 gnd vdd FILL
XFILL_47_DFFSR_73 gnd vdd FILL
XFILL_47_DFFSR_84 gnd vdd FILL
XFILL_61_DFFSR_242 gnd vdd FILL
XFILL_47_DFFSR_95 gnd vdd FILL
XFILL_61_DFFSR_253 gnd vdd FILL
XFILL_61_DFFSR_264 gnd vdd FILL
XFILL_61_DFFSR_275 gnd vdd FILL
XFILL_15_NOR3X1_30 gnd vdd FILL
XFILL_15_NOR3X1_41 gnd vdd FILL
XFILL_15_NOR3X1_52 gnd vdd FILL
XFILL_87_DFFSR_50 gnd vdd FILL
XFILL_87_DFFSR_61 gnd vdd FILL
XFILL_65_DFFSR_230 gnd vdd FILL
XFILL_87_DFFSR_72 gnd vdd FILL
XFILL_65_DFFSR_241 gnd vdd FILL
XFILL_87_DFFSR_83 gnd vdd FILL
XFILL_87_DFFSR_94 gnd vdd FILL
XFILL_65_DFFSR_252 gnd vdd FILL
XFILL_16_DFFSR_50 gnd vdd FILL
XFILL_16_DFFSR_61 gnd vdd FILL
XFILL_65_DFFSR_263 gnd vdd FILL
XFILL_65_DFFSR_274 gnd vdd FILL
XFILL_20_CLKBUF1_4 gnd vdd FILL
XFILL_16_DFFSR_72 gnd vdd FILL
XFILL_19_NOR3X1_40 gnd vdd FILL
XFILL_11_NAND2X1_19 gnd vdd FILL
XFILL_16_DFFSR_83 gnd vdd FILL
XFILL_19_NOR3X1_51 gnd vdd FILL
XFILL_60_2 gnd vdd FILL
XFILL_16_DFFSR_94 gnd vdd FILL
XFILL_27_NOR3X1_2 gnd vdd FILL
XFILL_69_DFFSR_240 gnd vdd FILL
XFILL_69_DFFSR_251 gnd vdd FILL
XFILL_53_1 gnd vdd FILL
XFILL_69_DFFSR_262 gnd vdd FILL
XFILL_56_DFFSR_60 gnd vdd FILL
XFILL_24_CLKBUF1_3 gnd vdd FILL
XFILL_69_DFFSR_273 gnd vdd FILL
XFILL_56_DFFSR_71 gnd vdd FILL
XFILL_56_DFFSR_82 gnd vdd FILL
XFILL_36_3_0 gnd vdd FILL
XFILL_2_NOR2X1_13 gnd vdd FILL
XFILL_56_DFFSR_93 gnd vdd FILL
XFILL_8_NAND3X1_12 gnd vdd FILL
XFILL_2_NOR2X1_24 gnd vdd FILL
XFILL_43_DFFSR_209 gnd vdd FILL
XFILL_8_NAND3X1_23 gnd vdd FILL
XFILL_2_NOR2X1_35 gnd vdd FILL
XFILL_8_NAND3X1_34 gnd vdd FILL
XFILL_2_NOR2X1_46 gnd vdd FILL
XFILL_1_NOR2X1_3 gnd vdd FILL
XFILL_8_NAND3X1_45 gnd vdd FILL
XFILL_2_NOR2X1_57 gnd vdd FILL
XFILL_8_NAND3X1_56 gnd vdd FILL
XFILL_2_NOR2X1_68 gnd vdd FILL
XFILL_28_CLKBUF1_2 gnd vdd FILL
XFILL_2_NOR2X1_79 gnd vdd FILL
XFILL_8_NAND3X1_67 gnd vdd FILL
XFILL_8_NAND3X1_78 gnd vdd FILL
XFILL_70_DFFSR_109 gnd vdd FILL
XFILL_8_NAND3X1_89 gnd vdd FILL
XFILL_6_NOR2X1_12 gnd vdd FILL
XFILL_47_DFFSR_208 gnd vdd FILL
XFILL_6_NOR2X1_23 gnd vdd FILL
XFILL_47_DFFSR_219 gnd vdd FILL
XFILL_9_OAI21X1_9 gnd vdd FILL
XFILL_25_DFFSR_70 gnd vdd FILL
XFILL_6_NOR2X1_34 gnd vdd FILL
XFILL_25_DFFSR_81 gnd vdd FILL
XFILL_6_NOR2X1_45 gnd vdd FILL
XFILL_6_NOR2X1_56 gnd vdd FILL
XFILL_25_DFFSR_92 gnd vdd FILL
XFILL_10_OAI22X1_7 gnd vdd FILL
XFILL_6_NOR2X1_67 gnd vdd FILL
XFILL_6_NOR2X1_78 gnd vdd FILL
XFILL_20_7_1 gnd vdd FILL
XFILL_0_MUX2X1_1 gnd vdd FILL
XFILL_6_NOR2X1_89 gnd vdd FILL
XFILL_74_DFFSR_108 gnd vdd FILL
XFILL_74_DFFSR_119 gnd vdd FILL
XFILL_65_DFFSR_80 gnd vdd FILL
XFILL_15_AOI21X1_19 gnd vdd FILL
XFILL_14_OAI22X1_6 gnd vdd FILL
XFILL_65_DFFSR_91 gnd vdd FILL
XFILL_1_NAND2X1_14 gnd vdd FILL
XFILL_6_DFFSR_3 gnd vdd FILL
XFILL_1_NAND2X1_25 gnd vdd FILL
XFILL_15_NAND3X1_110 gnd vdd FILL
XFILL_15_NAND3X1_121 gnd vdd FILL
XFILL_1_NAND2X1_36 gnd vdd FILL
XFILL_15_NAND3X1_132 gnd vdd FILL
XFILL_78_DFFSR_107 gnd vdd FILL
XFILL_19_DFFSR_1 gnd vdd FILL
XFILL_1_NAND2X1_47 gnd vdd FILL
XFILL_1_NAND2X1_58 gnd vdd FILL
XFILL_78_DFFSR_118 gnd vdd FILL
XFILL_1_NAND2X1_69 gnd vdd FILL
XFILL_76_DFFSR_2 gnd vdd FILL
XFILL_78_DFFSR_129 gnd vdd FILL
XFILL_8_DFFSR_60 gnd vdd FILL
XFILL_18_OAI22X1_5 gnd vdd FILL
XFILL_8_DFFSR_71 gnd vdd FILL
XFILL_8_DFFSR_82 gnd vdd FILL
XFILL_8_DFFSR_93 gnd vdd FILL
XFILL_34_DFFSR_90 gnd vdd FILL
XFILL_1_BUFX2_9 gnd vdd FILL
XFILL_32_DFFSR_230 gnd vdd FILL
XFILL_32_DFFSR_241 gnd vdd FILL
XFILL_6_NAND3X1_104 gnd vdd FILL
XFILL_6_NAND3X1_115 gnd vdd FILL
XFILL_32_DFFSR_252 gnd vdd FILL
XFILL_6_NAND3X1_126 gnd vdd FILL
XFILL_32_DFFSR_263 gnd vdd FILL
XFILL_32_DFFSR_274 gnd vdd FILL
XFILL_27_CLKBUF1_13 gnd vdd FILL
XFILL_27_CLKBUF1_24 gnd vdd FILL
XFILL_60_DFFSR_8 gnd vdd FILL
XFILL_27_CLKBUF1_35 gnd vdd FILL
XFILL_36_DFFSR_240 gnd vdd FILL
XFILL_27_3_0 gnd vdd FILL
XFILL_36_DFFSR_251 gnd vdd FILL
XFILL_2_3_0 gnd vdd FILL
XFILL_36_DFFSR_262 gnd vdd FILL
XFILL_36_DFFSR_273 gnd vdd FILL
XFILL_2_MUX2X1_20 gnd vdd FILL
XFILL_2_MUX2X1_31 gnd vdd FILL
XFILL_2_MUX2X1_42 gnd vdd FILL
XFILL_10_DFFSR_209 gnd vdd FILL
XFILL_2_MUX2X1_53 gnd vdd FILL
XFILL_5_AOI21X1_14 gnd vdd FILL
XFILL_2_MUX2X1_64 gnd vdd FILL
XFILL_5_AOI21X1_25 gnd vdd FILL
XFILL_63_DFFSR_140 gnd vdd FILL
XFILL_2_MUX2X1_75 gnd vdd FILL
XFILL_5_AOI21X1_36 gnd vdd FILL
XFILL_63_DFFSR_151 gnd vdd FILL
XFILL_63_DFFSR_162 gnd vdd FILL
XFILL_2_MUX2X1_86 gnd vdd FILL
XFILL_5_AOI21X1_47 gnd vdd FILL
XFILL_2_MUX2X1_97 gnd vdd FILL
XFILL_63_DFFSR_173 gnd vdd FILL
XFILL_15_OAI22X1_16 gnd vdd FILL
XFILL_5_AOI21X1_58 gnd vdd FILL
XFILL_5_AOI21X1_69 gnd vdd FILL
XFILL_63_DFFSR_184 gnd vdd FILL
XFILL_6_MUX2X1_30 gnd vdd FILL
XFILL_15_OAI22X1_27 gnd vdd FILL
XFILL_63_DFFSR_195 gnd vdd FILL
XFILL_15_OAI22X1_38 gnd vdd FILL
XFILL_14_DFFSR_208 gnd vdd FILL
XFILL_8_NOR2X1_102 gnd vdd FILL
XFILL_6_MUX2X1_41 gnd vdd FILL
XFILL_15_OAI22X1_49 gnd vdd FILL
XFILL_8_NOR2X1_113 gnd vdd FILL
XFILL_14_DFFSR_219 gnd vdd FILL
XFILL_6_MUX2X1_52 gnd vdd FILL
XFILL_11_NAND3X1_8 gnd vdd FILL
XFILL_8_NOR2X1_124 gnd vdd FILL
XFILL_11_7_1 gnd vdd FILL
XFILL_6_MUX2X1_63 gnd vdd FILL
XFILL_6_MUX2X1_74 gnd vdd FILL
XFILL_0_BUFX4_3 gnd vdd FILL
XFILL_67_DFFSR_150 gnd vdd FILL
XFILL_8_NOR2X1_135 gnd vdd FILL
XFILL_67_DFFSR_161 gnd vdd FILL
XFILL_8_NOR2X1_146 gnd vdd FILL
XFILL_6_MUX2X1_85 gnd vdd FILL
XFILL_10_2_0 gnd vdd FILL
XFILL_6_MUX2X1_96 gnd vdd FILL
XFILL_8_NOR2X1_157 gnd vdd FILL
XFILL_67_DFFSR_172 gnd vdd FILL
XFILL_13_BUFX4_1 gnd vdd FILL
XFILL_67_DFFSR_183 gnd vdd FILL
XFILL_8_NOR2X1_168 gnd vdd FILL
XFILL_8_NOR2X1_179 gnd vdd FILL
XFILL_41_DFFSR_108 gnd vdd FILL
XFILL_67_DFFSR_194 gnd vdd FILL
XFILL_18_DFFSR_207 gnd vdd FILL
XFILL_14_NAND3X1_70 gnd vdd FILL
XFILL_15_NAND3X1_7 gnd vdd FILL
XFILL_14_NAND3X1_81 gnd vdd FILL
XFILL_41_DFFSR_119 gnd vdd FILL
XFILL_18_DFFSR_218 gnd vdd FILL
XFILL_14_NAND3X1_92 gnd vdd FILL
XFILL_18_DFFSR_229 gnd vdd FILL
XFILL_1_NAND3X1_100 gnd vdd FILL
XFILL_1_NAND3X1_111 gnd vdd FILL
XFILL_1_NAND3X1_122 gnd vdd FILL
XFILL_45_DFFSR_107 gnd vdd FILL
XFILL_45_DFFSR_118 gnd vdd FILL
XFILL_45_DFFSR_129 gnd vdd FILL
XFILL_49_DFFSR_106 gnd vdd FILL
XFILL_8_MUX2X1_108 gnd vdd FILL
XFILL_8_MUX2X1_119 gnd vdd FILL
XFILL_49_DFFSR_117 gnd vdd FILL
XFILL_49_DFFSR_128 gnd vdd FILL
XFILL_49_DFFSR_139 gnd vdd FILL
XFILL_22_MUX2X1_50 gnd vdd FILL
XFILL_5_OAI22X1_11 gnd vdd FILL
XFILL_22_MUX2X1_61 gnd vdd FILL
XFILL_11_AND2X2_8 gnd vdd FILL
XFILL_5_OAI22X1_22 gnd vdd FILL
XFILL_22_MUX2X1_72 gnd vdd FILL
XFILL_5_OAI22X1_33 gnd vdd FILL
XFILL_22_MUX2X1_83 gnd vdd FILL
XFILL_5_OAI22X1_44 gnd vdd FILL
XFILL_22_MUX2X1_94 gnd vdd FILL
XFILL_9_OAI21X1_13 gnd vdd FILL
XFILL_9_OAI21X1_24 gnd vdd FILL
XFILL_18_3_0 gnd vdd FILL
XFILL_9_OAI21X1_35 gnd vdd FILL
XFILL_9_OAI21X1_46 gnd vdd FILL
XFILL_32_6 gnd vdd FILL
XFILL_61_6_1 gnd vdd FILL
XFILL_60_1_0 gnd vdd FILL
XFILL_25_5 gnd vdd FILL
XFILL_2_NOR2X1_202 gnd vdd FILL
XFILL_30_DFFSR_140 gnd vdd FILL
XFILL_3_INVX8_1 gnd vdd FILL
XFILL_30_DFFSR_151 gnd vdd FILL
XFILL_30_DFFSR_162 gnd vdd FILL
XFILL_18_4 gnd vdd FILL
XFILL_30_DFFSR_173 gnd vdd FILL
XFILL_30_DFFSR_184 gnd vdd FILL
XFILL_30_DFFSR_195 gnd vdd FILL
XFILL_16_CLKBUF1_20 gnd vdd FILL
XFILL_16_CLKBUF1_31 gnd vdd FILL
XFILL_16_CLKBUF1_42 gnd vdd FILL
XFILL_34_DFFSR_150 gnd vdd FILL
XFILL_34_DFFSR_161 gnd vdd FILL
XFILL_34_DFFSR_172 gnd vdd FILL
XFILL_11_AOI21X1_50 gnd vdd FILL
XFILL_34_DFFSR_183 gnd vdd FILL
XFILL_79_DFFSR_19 gnd vdd FILL
XFILL_34_DFFSR_194 gnd vdd FILL
XFILL_20_DFFSR_1 gnd vdd FILL
XFILL_11_AOI21X1_61 gnd vdd FILL
XFILL_11_AOI21X1_72 gnd vdd FILL
XFILL_38_DFFSR_160 gnd vdd FILL
XFILL_2_INVX1_15 gnd vdd FILL
XFILL_38_DFFSR_171 gnd vdd FILL
XFILL_2_INVX1_26 gnd vdd FILL
XFILL_38_DFFSR_182 gnd vdd FILL
XFILL_12_DFFSR_107 gnd vdd FILL
XFILL_2_INVX1_37 gnd vdd FILL
XFILL_38_DFFSR_193 gnd vdd FILL
XFILL_2_INVX1_48 gnd vdd FILL
XFILL_3_AND2X2_7 gnd vdd FILL
XFILL_30_NOR3X1_40 gnd vdd FILL
XFILL_2_INVX1_59 gnd vdd FILL
XFILL_12_DFFSR_118 gnd vdd FILL
XFILL_30_NOR3X1_51 gnd vdd FILL
XFILL_12_DFFSR_129 gnd vdd FILL
XFILL_48_DFFSR_18 gnd vdd FILL
XFILL_48_DFFSR_29 gnd vdd FILL
XFILL_80_DFFSR_240 gnd vdd FILL
XFILL_80_DFFSR_251 gnd vdd FILL
XFILL_80_DFFSR_262 gnd vdd FILL
XFILL_16_DFFSR_106 gnd vdd FILL
XFILL_80_DFFSR_273 gnd vdd FILL
XFILL_16_DFFSR_117 gnd vdd FILL
XFILL_16_DFFSR_128 gnd vdd FILL
XFILL_16_DFFSR_139 gnd vdd FILL
XFILL_0_BUFX4_13 gnd vdd FILL
XFILL_11_AOI21X1_2 gnd vdd FILL
XFILL_42_DFFSR_5 gnd vdd FILL
XFILL_0_BUFX4_24 gnd vdd FILL
XFILL_0_BUFX4_35 gnd vdd FILL
XFILL_84_DFFSR_250 gnd vdd FILL
XFILL_0_BUFX4_46 gnd vdd FILL
XFILL_84_DFFSR_261 gnd vdd FILL
XFILL_0_BUFX4_57 gnd vdd FILL
XFILL_84_DFFSR_272 gnd vdd FILL
XFILL_17_DFFSR_17 gnd vdd FILL
XFILL_0_BUFX4_68 gnd vdd FILL
XFILL_17_DFFSR_28 gnd vdd FILL
XFILL_14_MUX2X1_100 gnd vdd FILL
XFILL_17_DFFSR_39 gnd vdd FILL
XFILL_14_MUX2X1_111 gnd vdd FILL
XFILL_0_BUFX4_79 gnd vdd FILL
XFILL_14_MUX2X1_122 gnd vdd FILL
XFILL_52_6_1 gnd vdd FILL
XFILL_15_AOI21X1_1 gnd vdd FILL
XFILL_14_MUX2X1_133 gnd vdd FILL
XFILL_14_MUX2X1_144 gnd vdd FILL
XFILL_51_1_0 gnd vdd FILL
XFILL_14_MUX2X1_155 gnd vdd FILL
XFILL_12_NOR3X1_18 gnd vdd FILL
XFILL_57_DFFSR_16 gnd vdd FILL
XFILL_14_MUX2X1_166 gnd vdd FILL
XFILL_12_NOR3X1_29 gnd vdd FILL
XFILL_14_MUX2X1_177 gnd vdd FILL
XFILL_57_DFFSR_27 gnd vdd FILL
XFILL_14_MUX2X1_188 gnd vdd FILL
XFILL_57_DFFSR_38 gnd vdd FILL
XFILL_62_DFFSR_207 gnd vdd FILL
XFILL_57_DFFSR_49 gnd vdd FILL
XFILL_62_DFFSR_218 gnd vdd FILL
XFILL_62_DFFSR_229 gnd vdd FILL
XFILL_16_NOR3X1_17 gnd vdd FILL
XFILL_16_NOR3X1_28 gnd vdd FILL
XFILL_16_NOR3X1_39 gnd vdd FILL
XFILL_66_DFFSR_206 gnd vdd FILL
XFILL_64_DFFSR_9 gnd vdd FILL
XFILL_66_DFFSR_217 gnd vdd FILL
XFILL_26_DFFSR_15 gnd vdd FILL
XFILL_26_DFFSR_26 gnd vdd FILL
XFILL_66_DFFSR_228 gnd vdd FILL
XFILL_66_DFFSR_239 gnd vdd FILL
XFILL_26_DFFSR_37 gnd vdd FILL
XFILL_26_DFFSR_48 gnd vdd FILL
XFILL_26_DFFSR_59 gnd vdd FILL
XFILL_66_DFFSR_14 gnd vdd FILL
XFILL_66_DFFSR_25 gnd vdd FILL
XFILL_66_DFFSR_36 gnd vdd FILL
XFILL_66_DFFSR_47 gnd vdd FILL
XFILL_66_DFFSR_58 gnd vdd FILL
XFILL_66_DFFSR_69 gnd vdd FILL
XNAND3X1_13 DFFSR_1/D NAND3X1_43/B OAI21X1_42/Y gnd NOR3X1_52/C vdd NAND3X1
XFILL_59_2_0 gnd vdd FILL
XFILL_21_MUX2X1_190 gnd vdd FILL
XNAND3X1_24 NAND3X1_67/Y OAI21X1_23/Y NOR3X1_9/A gnd NOR2X1_37/B vdd NAND3X1
XNAND3X1_35 NAND3X1_43/A NAND3X1_39/B OAI21X1_45/Y gnd NOR3X1_2/C vdd NAND3X1
XFILL_4_MUX2X1_150 gnd vdd FILL
XNAND3X1_46 NAND3X1_46/A NAND3X1_46/B NAND3X1_46/C gnd NOR2X1_39/B vdd NAND3X1
XFILL_4_BUFX4_4 gnd vdd FILL
XNAND3X1_57 AND2X2_1/B AND2X2_6/A BUFX4_57/Y gnd OAI22X1_7/B vdd NAND3X1
XFILL_9_DFFSR_16 gnd vdd FILL
XFILL_4_MUX2X1_161 gnd vdd FILL
XFILL_9_DFFSR_27 gnd vdd FILL
XNAND3X1_68 INVX2_2/A OAI21X1_50/Y NOR2X1_54/Y gnd NOR3X1_46/B vdd NAND3X1
XFILL_4_MUX2X1_172 gnd vdd FILL
XFILL_7_NAND3X1_105 gnd vdd FILL
XFILL_35_DFFSR_13 gnd vdd FILL
XFILL_9_DFFSR_38 gnd vdd FILL
XFILL_7_NAND3X1_116 gnd vdd FILL
XNAND3X1_79 DFFSR_20/Q NAND3X1_7/B NOR2X1_34/Y gnd NAND3X1_82/A vdd NAND3X1
XFILL_4_MUX2X1_183 gnd vdd FILL
XFILL_35_DFFSR_24 gnd vdd FILL
XFILL_4_MUX2X1_194 gnd vdd FILL
XFILL_9_DFFSR_49 gnd vdd FILL
XFILL_7_NAND3X1_127 gnd vdd FILL
XFILL_35_DFFSR_35 gnd vdd FILL
XNOR2X1_13 INVX2_3/A NOR2X1_13/B gnd NOR2X1_13/Y vdd NOR2X1
XFILL_35_DFFSR_46 gnd vdd FILL
XNOR2X1_24 NOR2X1_24/A NOR2X1_24/B gnd NOR2X1_24/Y vdd NOR2X1
XNOR2X1_35 INVX4_1/Y NOR2X1_35/B gnd NOR2X1_46/B vdd NOR2X1
XFILL_35_DFFSR_57 gnd vdd FILL
XNOR2X1_46 NOR2X1_46/A NOR2X1_46/B gnd NOR2X1_46/Y vdd NOR2X1
XFILL_35_DFFSR_68 gnd vdd FILL
XFILL_35_DFFSR_79 gnd vdd FILL
XNOR2X1_57 NOR2X1_57/A INVX4_1/Y gnd NOR2X1_57/Y vdd NOR2X1
XNOR2X1_68 NOR2X1_68/A INVX4_1/Y gnd NOR2X1_90/B vdd NOR2X1
XNOR2X1_79 NOR2X1_79/A NOR2X1_90/B gnd NOR2X1_79/Y vdd NOR2X1
XFILL_75_DFFSR_12 gnd vdd FILL
XFILL_51_DFFSR_250 gnd vdd FILL
XFILL_75_DFFSR_23 gnd vdd FILL
XFILL_51_DFFSR_261 gnd vdd FILL
XFILL_43_6_1 gnd vdd FILL
XFILL_51_DFFSR_272 gnd vdd FILL
XFILL_75_DFFSR_34 gnd vdd FILL
XFILL_75_DFFSR_45 gnd vdd FILL
XFILL_75_DFFSR_56 gnd vdd FILL
XFILL_18_MUX2X1_2 gnd vdd FILL
XFILL_42_1_0 gnd vdd FILL
XFILL_75_DFFSR_67 gnd vdd FILL
XFILL_75_DFFSR_78 gnd vdd FILL
XFILL_75_DFFSR_89 gnd vdd FILL
XFILL_3_INVX1_8 gnd vdd FILL
XFILL_55_DFFSR_260 gnd vdd FILL
XFILL_55_DFFSR_271 gnd vdd FILL
XFILL_10_CLKBUF1_1 gnd vdd FILL
XFILL_10_NAND2X1_16 gnd vdd FILL
XFILL_10_NAND2X1_27 gnd vdd FILL
XFILL_44_DFFSR_11 gnd vdd FILL
XFILL_10_NAND2X1_38 gnd vdd FILL
XFILL_10_NAND2X1_49 gnd vdd FILL
XFILL_44_DFFSR_22 gnd vdd FILL
XFILL_44_DFFSR_33 gnd vdd FILL
XFILL_15_NOR3X1_8 gnd vdd FILL
XFILL_9_BUFX4_90 gnd vdd FILL
XFILL_44_DFFSR_44 gnd vdd FILL
XFILL_44_DFFSR_55 gnd vdd FILL
XFILL_82_DFFSR_160 gnd vdd FILL
XFILL_44_DFFSR_66 gnd vdd FILL
XFILL_82_DFFSR_171 gnd vdd FILL
XFILL_44_DFFSR_77 gnd vdd FILL
XFILL_59_DFFSR_270 gnd vdd FILL
XFILL_44_DFFSR_88 gnd vdd FILL
XFILL_82_DFFSR_182 gnd vdd FILL
XFILL_44_DFFSR_99 gnd vdd FILL
XFILL_82_DFFSR_193 gnd vdd FILL
XFILL_84_DFFSR_10 gnd vdd FILL
XFILL_33_DFFSR_206 gnd vdd FILL
XFILL_84_DFFSR_21 gnd vdd FILL
XFILL_7_NAND3X1_20 gnd vdd FILL
XFILL_33_DFFSR_217 gnd vdd FILL
XFILL_2_DFFSR_230 gnd vdd FILL
XFILL_2_DFFSR_241 gnd vdd FILL
XFILL_33_DFFSR_228 gnd vdd FILL
XFILL_84_DFFSR_32 gnd vdd FILL
XFILL_84_DFFSR_43 gnd vdd FILL
XFILL_2_NAND3X1_101 gnd vdd FILL
XFILL_7_NAND3X1_31 gnd vdd FILL
XFILL_33_DFFSR_239 gnd vdd FILL
XFILL_2_DFFSR_252 gnd vdd FILL
XFILL_13_DFFSR_10 gnd vdd FILL
XFILL_84_DFFSR_54 gnd vdd FILL
XFILL_7_NAND3X1_42 gnd vdd FILL
XFILL_2_NAND3X1_112 gnd vdd FILL
XFILL_13_DFFSR_21 gnd vdd FILL
XFILL_84_DFFSR_65 gnd vdd FILL
XFILL_7_NAND3X1_53 gnd vdd FILL
XFILL_2_NAND3X1_123 gnd vdd FILL
XFILL_2_DFFSR_263 gnd vdd FILL
XFILL_84_DFFSR_76 gnd vdd FILL
XFILL_2_DFFSR_274 gnd vdd FILL
XFILL_86_DFFSR_170 gnd vdd FILL
XFILL_7_NAND3X1_64 gnd vdd FILL
XFILL_13_DFFSR_32 gnd vdd FILL
XFILL_86_DFFSR_181 gnd vdd FILL
XFILL_13_DFFSR_43 gnd vdd FILL
XFILL_7_NAND3X1_75 gnd vdd FILL
XFILL_84_DFFSR_87 gnd vdd FILL
XFILL_60_DFFSR_106 gnd vdd FILL
XFILL_84_DFFSR_98 gnd vdd FILL
XFILL_7_NAND3X1_86 gnd vdd FILL
XFILL_86_DFFSR_192 gnd vdd FILL
XFILL_13_DFFSR_54 gnd vdd FILL
XFILL_37_DFFSR_205 gnd vdd FILL
XFILL_7_NAND3X1_97 gnd vdd FILL
XFILL_13_DFFSR_65 gnd vdd FILL
XFILL_60_DFFSR_117 gnd vdd FILL
XFILL_13_DFFSR_76 gnd vdd FILL
XFILL_37_DFFSR_216 gnd vdd FILL
XFILL_37_DFFSR_227 gnd vdd FILL
XFILL_6_DFFSR_240 gnd vdd FILL
XFILL_60_DFFSR_128 gnd vdd FILL
XFILL_7_INVX8_2 gnd vdd FILL
XFILL_6_DFFSR_251 gnd vdd FILL
XFILL_37_DFFSR_238 gnd vdd FILL
XFILL_13_DFFSR_87 gnd vdd FILL
XFILL_60_DFFSR_139 gnd vdd FILL
XFILL_13_DFFSR_98 gnd vdd FILL
XFILL_37_DFFSR_249 gnd vdd FILL
XFILL_6_DFFSR_262 gnd vdd FILL
XFILL_53_DFFSR_20 gnd vdd FILL
XFILL_6_DFFSR_273 gnd vdd FILL
XFILL_53_DFFSR_31 gnd vdd FILL
XFILL_3_MUX2X1_18 gnd vdd FILL
XFILL_24_NOR3X1_6 gnd vdd FILL
XFILL_53_DFFSR_42 gnd vdd FILL
XFILL_64_DFFSR_105 gnd vdd FILL
XFILL_3_MUX2X1_29 gnd vdd FILL
XFILL_53_DFFSR_53 gnd vdd FILL
XFILL_19_CLKBUF1_19 gnd vdd FILL
XFILL_64_DFFSR_116 gnd vdd FILL
XFILL_53_DFFSR_64 gnd vdd FILL
XFILL_53_DFFSR_75 gnd vdd FILL
XFILL_53_DFFSR_86 gnd vdd FILL
XFILL_64_DFFSR_127 gnd vdd FILL
XFILL_64_DFFSR_138 gnd vdd FILL
XFILL_64_DFFSR_149 gnd vdd FILL
XFILL_14_AOI21X1_16 gnd vdd FILL
XFILL_53_DFFSR_97 gnd vdd FILL
XFILL_0_NAND2X1_11 gnd vdd FILL
XFILL_14_AOI21X1_27 gnd vdd FILL
XFILL_0_NAND2X1_22 gnd vdd FILL
XMUX2X1_20 BUFX4_97/Y INVX1_33/Y MUX2X1_20/S gnd DFFSR_14/D vdd MUX2X1
XMUX2X1_31 BUFX4_71/Y INVX1_44/Y NOR2X1_19/B gnd MUX2X1_31/Y vdd MUX2X1
XFILL_14_AOI21X1_38 gnd vdd FILL
XFILL_7_MUX2X1_17 gnd vdd FILL
XFILL_0_NAND2X1_33 gnd vdd FILL
XFILL_14_AOI21X1_49 gnd vdd FILL
XNOR2X1_103 OAI22X1_42/Y OAI22X1_43/Y gnd NOR2X1_103/Y vdd NOR2X1
XFILL_0_NAND2X1_44 gnd vdd FILL
XMUX2X1_42 INVX1_55/Y MUX2X1_9/A NAND2X1_6/Y gnd MUX2X1_42/Y vdd MUX2X1
XFILL_24_DFFSR_2 gnd vdd FILL
XFILL_7_MUX2X1_28 gnd vdd FILL
XFILL_68_DFFSR_104 gnd vdd FILL
XNOR2X1_114 INVX1_132/A INVX1_130/Y gnd OAI21X1_1/B vdd NOR2X1
XFILL_81_DFFSR_3 gnd vdd FILL
XFILL_0_NAND2X1_55 gnd vdd FILL
XMUX2X1_53 INVX1_66/Y MUX2X1_66/A NAND2X1_8/Y gnd MUX2X1_53/Y vdd MUX2X1
XFILL_7_MUX2X1_39 gnd vdd FILL
XFILL_68_DFFSR_115 gnd vdd FILL
XNOR2X1_125 DFFSR_149/Q AOI21X1_3/B gnd NOR2X1_125/Y vdd NOR2X1
XFILL_0_NAND2X1_66 gnd vdd FILL
XMUX2X1_64 BUFX4_63/Y INVX1_77/Y NOR2X1_23/Y gnd MUX2X1_64/Y vdd MUX2X1
XFILL_68_DFFSR_126 gnd vdd FILL
XFILL_22_DFFSR_30 gnd vdd FILL
XMUX2X1_75 INVX1_88/Y BUFX4_96/Y OR2X2_1/Y gnd MUX2X1_75/Y vdd MUX2X1
XFILL_0_NAND2X1_77 gnd vdd FILL
XFILL_22_DFFSR_41 gnd vdd FILL
XNOR2X1_136 INVX4_1/Y NOR2X1_10/B gnd NOR2X1_136/Y vdd NOR2X1
XFILL_68_DFFSR_137 gnd vdd FILL
XNOR2X1_147 DFFSR_106/Q AOI21X1_9/B gnd NOR2X1_147/Y vdd NOR2X1
XMUX2X1_86 INVX1_99/Y BUFX4_96/Y MUX2X1_86/S gnd MUX2X1_86/Y vdd MUX2X1
XFILL_34_6_1 gnd vdd FILL
XFILL_0_NAND2X1_88 gnd vdd FILL
XFILL_68_DFFSR_148 gnd vdd FILL
XFILL_11_OAI21X1_5 gnd vdd FILL
XMUX2X1_97 NOR2X1_60/A BUFX4_64/Y MUX2X1_99/S gnd DFFSR_68/D vdd MUX2X1
XNOR2X1_158 DFFSR_81/Q NOR2X1_161/B gnd NOR2X1_158/Y vdd NOR2X1
XFILL_22_DFFSR_52 gnd vdd FILL
XFILL_22_DFFSR_63 gnd vdd FILL
XFILL_68_DFFSR_159 gnd vdd FILL
XNOR2X1_169 NAND2X1_3/Y INVX1_8/Y gnd NOR2X1_169/Y vdd NOR2X1
XFILL_22_DFFSR_74 gnd vdd FILL
XFILL_33_1_0 gnd vdd FILL
XFILL_22_DFFSR_85 gnd vdd FILL
XFILL_22_DFFSR_96 gnd vdd FILL
XFILL_23_2 gnd vdd FILL
XFILL_7_NOR3X1_7 gnd vdd FILL
XFILL_62_DFFSR_40 gnd vdd FILL
XFILL_62_DFFSR_51 gnd vdd FILL
XFILL_3_AOI22X1_1 gnd vdd FILL
XFILL_16_1 gnd vdd FILL
XFILL_15_OAI21X1_4 gnd vdd FILL
XFILL_62_DFFSR_62 gnd vdd FILL
XFILL_62_DFFSR_73 gnd vdd FILL
XFILL_62_DFFSR_84 gnd vdd FILL
XFILL_22_DFFSR_260 gnd vdd FILL
XFILL_62_DFFSR_95 gnd vdd FILL
XFILL_22_DFFSR_271 gnd vdd FILL
XFILL_3_INVX1_200 gnd vdd FILL
XFILL_26_CLKBUF1_10 gnd vdd FILL
XFILL_3_INVX1_211 gnd vdd FILL
XFILL_26_CLKBUF1_21 gnd vdd FILL
XDFFSR_1 INVX2_4/A DFFSR_1/CLK DFFSR_1/R vdd DFFSR_1/D gnd vdd DFFSR
XFILL_3_INVX1_222 gnd vdd FILL
XFILL_26_CLKBUF1_32 gnd vdd FILL
XFILL_5_DFFSR_20 gnd vdd FILL
XFILL_5_DFFSR_31 gnd vdd FILL
XFILL_5_DFFSR_42 gnd vdd FILL
XFILL_46_DFFSR_6 gnd vdd FILL
XFILL_5_DFFSR_53 gnd vdd FILL
XMUX2X1_109 NOR2X1_47/A BUFX4_80/Y NAND2X1_23/Y gnd DFFSR_152/D vdd MUX2X1
XFILL_5_DFFSR_64 gnd vdd FILL
XFILL_26_DFFSR_270 gnd vdd FILL
XFILL_5_DFFSR_75 gnd vdd FILL
XFILL_9_CLKBUF1_14 gnd vdd FILL
XFILL_31_DFFSR_50 gnd vdd FILL
XFILL_9_CLKBUF1_25 gnd vdd FILL
XFILL_5_DFFSR_86 gnd vdd FILL
XFILL_23_MUX2X1_15 gnd vdd FILL
XFILL_31_DFFSR_61 gnd vdd FILL
XFILL_7_INVX1_210 gnd vdd FILL
XFILL_9_CLKBUF1_36 gnd vdd FILL
XFILL_23_MUX2X1_26 gnd vdd FILL
XFILL_5_DFFSR_97 gnd vdd FILL
XFILL_7_INVX1_221 gnd vdd FILL
XFILL_31_DFFSR_72 gnd vdd FILL
XFILL_31_DFFSR_83 gnd vdd FILL
XFILL_4_AOI21X1_11 gnd vdd FILL
XFILL_23_MUX2X1_37 gnd vdd FILL
XFILL_4_AOI21X1_22 gnd vdd FILL
XFILL_23_MUX2X1_48 gnd vdd FILL
XFILL_31_DFFSR_94 gnd vdd FILL
XFILL_4_AOI21X1_33 gnd vdd FILL
XFILL_23_MUX2X1_59 gnd vdd FILL
XFILL_4_AOI21X1_44 gnd vdd FILL
XFILL_53_DFFSR_170 gnd vdd FILL
XFILL_4_AOI21X1_55 gnd vdd FILL
XFILL_14_OAI22X1_13 gnd vdd FILL
XFILL_4_AOI21X1_66 gnd vdd FILL
XFILL_14_OAI22X1_24 gnd vdd FILL
XFILL_53_DFFSR_181 gnd vdd FILL
XFILL_4_AOI21X1_77 gnd vdd FILL
XFILL_71_DFFSR_60 gnd vdd FILL
XFILL_14_OAI22X1_35 gnd vdd FILL
XFILL_53_DFFSR_192 gnd vdd FILL
XFILL_71_DFFSR_71 gnd vdd FILL
XFILL_14_OAI22X1_46 gnd vdd FILL
XINVX1_16 INVX1_16/A gnd MUX2X1_3/B vdd INVX1
XFILL_71_DFFSR_82 gnd vdd FILL
XFILL_7_NOR2X1_110 gnd vdd FILL
XINVX1_27 INVX1_27/A gnd INVX1_27/Y vdd INVX1
XINVX1_38 INVX1_38/A gnd INVX1_38/Y vdd INVX1
XFILL_71_DFFSR_93 gnd vdd FILL
XFILL_7_NOR2X1_121 gnd vdd FILL
XFILL_7_NOR2X1_132 gnd vdd FILL
XINVX1_49 INVX1_49/A gnd INVX1_49/Y vdd INVX1
XFILL_7_NOR2X1_143 gnd vdd FILL
XFILL_7_NOR2X1_154 gnd vdd FILL
XFILL_57_DFFSR_180 gnd vdd FILL
XFILL_7_NOR2X1_165 gnd vdd FILL
XFILL_7_NOR2X1_176 gnd vdd FILL
XFILL_7_NOR2X1_187 gnd vdd FILL
XFILL_31_DFFSR_105 gnd vdd FILL
XFILL_57_DFFSR_191 gnd vdd FILL
XFILL_31_DFFSR_116 gnd vdd FILL
XFILL_11_NOR3X1_1 gnd vdd FILL
XFILL_7_NOR2X1_198 gnd vdd FILL
XFILL_0_DFFSR_140 gnd vdd FILL
XFILL_31_DFFSR_127 gnd vdd FILL
XNAND2X1_90 INVX1_139/A NOR2X1_21/B gnd NAND3X1_30/C vdd NAND2X1
XFILL_31_DFFSR_138 gnd vdd FILL
XFILL_0_DFFSR_151 gnd vdd FILL
XFILL_11_NOR2X1_204 gnd vdd FILL
XFILL_0_DFFSR_162 gnd vdd FILL
XFILL_31_DFFSR_149 gnd vdd FILL
XFILL_40_DFFSR_70 gnd vdd FILL
XFILL_0_DFFSR_173 gnd vdd FILL
XFILL_40_DFFSR_81 gnd vdd FILL
XFILL_0_DFFSR_184 gnd vdd FILL
XFILL_40_DFFSR_92 gnd vdd FILL
XFILL_25_6_1 gnd vdd FILL
XFILL_0_DFFSR_195 gnd vdd FILL
XFILL_35_DFFSR_104 gnd vdd FILL
XFILL_0_6_1 gnd vdd FILL
XFILL_35_DFFSR_115 gnd vdd FILL
XFILL_35_DFFSR_126 gnd vdd FILL
XFILL_24_1_0 gnd vdd FILL
XFILL_35_DFFSR_137 gnd vdd FILL
XFILL_4_DFFSR_150 gnd vdd FILL
XFILL_4_DFFSR_161 gnd vdd FILL
XFILL_35_DFFSR_148 gnd vdd FILL
XFILL_80_DFFSR_80 gnd vdd FILL
XFILL_4_DFFSR_172 gnd vdd FILL
XFILL_35_DFFSR_159 gnd vdd FILL
XFILL_4_DFFSR_183 gnd vdd FILL
XFILL_80_DFFSR_91 gnd vdd FILL
XFILL_4_DFFSR_194 gnd vdd FILL
XFILL_39_DFFSR_103 gnd vdd FILL
XFILL_7_MUX2X1_105 gnd vdd FILL
XFILL_7_MUX2X1_116 gnd vdd FILL
XFILL_39_DFFSR_114 gnd vdd FILL
XFILL_7_MUX2X1_127 gnd vdd FILL
XFILL_39_DFFSR_125 gnd vdd FILL
XFILL_39_DFFSR_136 gnd vdd FILL
XFILL_7_MUX2X1_138 gnd vdd FILL
XFILL_7_MUX2X1_149 gnd vdd FILL
XFILL_8_BUFX4_5 gnd vdd FILL
XFILL_8_DFFSR_160 gnd vdd FILL
XFILL_39_DFFSR_147 gnd vdd FILL
XFILL_39_DFFSR_158 gnd vdd FILL
XFILL_8_DFFSR_171 gnd vdd FILL
XFILL_12_MUX2X1_80 gnd vdd FILL
XFILL_4_OAI22X1_30 gnd vdd FILL
XFILL_39_DFFSR_169 gnd vdd FILL
XFILL_8_DFFSR_182 gnd vdd FILL
XFILL_4_OAI22X1_41 gnd vdd FILL
XFILL_31_NOR3X1_16 gnd vdd FILL
XFILL_12_MUX2X1_91 gnd vdd FILL
XFILL_8_DFFSR_193 gnd vdd FILL
XFILL_31_NOR3X1_27 gnd vdd FILL
XFILL_8_OAI21X1_10 gnd vdd FILL
XFILL_0_NOR3X1_40 gnd vdd FILL
XFILL_0_NOR3X1_51 gnd vdd FILL
XFILL_8_OAI21X1_21 gnd vdd FILL
XFILL_31_NOR3X1_38 gnd vdd FILL
XFILL_31_NOR3X1_49 gnd vdd FILL
XFILL_81_DFFSR_205 gnd vdd FILL
XFILL_8_OAI21X1_32 gnd vdd FILL
XFILL_81_DFFSR_216 gnd vdd FILL
XFILL_8_OAI21X1_43 gnd vdd FILL
XFILL_81_DFFSR_227 gnd vdd FILL
XFILL_81_DFFSR_238 gnd vdd FILL
XFILL_16_MUX2X1_90 gnd vdd FILL
XFILL_81_DFFSR_249 gnd vdd FILL
XFILL_4_NOR3X1_50 gnd vdd FILL
XFILL_85_DFFSR_204 gnd vdd FILL
XFILL_85_DFFSR_215 gnd vdd FILL
XFILL_85_DFFSR_226 gnd vdd FILL
XFILL_85_DFFSR_237 gnd vdd FILL
XFILL_8_7_1 gnd vdd FILL
XFILL_7_INVX1_9 gnd vdd FILL
XFILL_85_DFFSR_248 gnd vdd FILL
XFILL_20_DFFSR_170 gnd vdd FILL
XFILL_7_2_0 gnd vdd FILL
XFILL_85_DFFSR_259 gnd vdd FILL
XFILL_1_INVX1_110 gnd vdd FILL
XFILL_20_DFFSR_181 gnd vdd FILL
XFILL_1_INVX1_121 gnd vdd FILL
XFILL_20_DFFSR_192 gnd vdd FILL
XFILL_4_BUFX2_1 gnd vdd FILL
XFILL_1_INVX1_132 gnd vdd FILL
XFILL_1_INVX1_143 gnd vdd FILL
XFILL_1_INVX1_154 gnd vdd FILL
XFILL_1_INVX1_165 gnd vdd FILL
XFILL_1_INVX1_176 gnd vdd FILL
XFILL_8_NAND3X1_106 gnd vdd FILL
XFILL_24_DFFSR_180 gnd vdd FILL
XFILL_8_NAND3X1_117 gnd vdd FILL
XFILL_1_INVX1_187 gnd vdd FILL
XFILL_8_NAND3X1_128 gnd vdd FILL
XFILL_1_INVX1_198 gnd vdd FILL
XFILL_5_INVX1_120 gnd vdd FILL
XFILL_24_DFFSR_191 gnd vdd FILL
XFILL_5_INVX1_131 gnd vdd FILL
XFILL_10_AOI21X1_80 gnd vdd FILL
XFILL_5_INVX1_142 gnd vdd FILL
XFILL_5_INVX1_153 gnd vdd FILL
XFILL_5_INVX1_164 gnd vdd FILL
XFILL_16_6_1 gnd vdd FILL
XFILL_5_INVX1_175 gnd vdd FILL
XFILL_15_1_0 gnd vdd FILL
XFILL_1_DFFSR_90 gnd vdd FILL
XFILL_5_INVX1_186 gnd vdd FILL
XFILL_5_INVX1_197 gnd vdd FILL
XFILL_28_DFFSR_190 gnd vdd FILL
XFILL_12_NAND3X1_130 gnd vdd FILL
XFILL_70_DFFSR_270 gnd vdd FILL
XFILL_3_OAI22X1_4 gnd vdd FILL
XFILL_28_DFFSR_3 gnd vdd FILL
XFILL_85_DFFSR_4 gnd vdd FILL
XFILL_7_OAI22X1_3 gnd vdd FILL
XFILL_13_MUX2X1_130 gnd vdd FILL
XFILL_4_INVX2_1 gnd vdd FILL
XFILL_3_NAND3X1_102 gnd vdd FILL
XFILL_3_NAND3X1_113 gnd vdd FILL
XFILL_13_MUX2X1_141 gnd vdd FILL
XFILL_3_NAND3X1_124 gnd vdd FILL
XFILL_13_MUX2X1_152 gnd vdd FILL
XFILL_13_MUX2X1_163 gnd vdd FILL
XFILL_13_MUX2X1_174 gnd vdd FILL
XFILL_13_MUX2X1_185 gnd vdd FILL
XFILL_52_DFFSR_204 gnd vdd FILL
XFILL_52_DFFSR_215 gnd vdd FILL
XFILL_52_DFFSR_226 gnd vdd FILL
XFILL_52_DFFSR_237 gnd vdd FILL
XFILL_52_DFFSR_248 gnd vdd FILL
XFILL_52_DFFSR_259 gnd vdd FILL
XFILL_66_5_1 gnd vdd FILL
XFILL_12_DFFSR_9 gnd vdd FILL
XFILL_56_DFFSR_203 gnd vdd FILL
XFILL_65_0_0 gnd vdd FILL
XFILL_56_DFFSR_214 gnd vdd FILL
XFILL_56_DFFSR_225 gnd vdd FILL
XFILL_56_DFFSR_236 gnd vdd FILL
XFILL_56_DFFSR_247 gnd vdd FILL
XFILL_56_DFFSR_258 gnd vdd FILL
XFILL_56_DFFSR_269 gnd vdd FILL
XFILL_83_DFFSR_103 gnd vdd FILL
XFILL_83_DFFSR_114 gnd vdd FILL
XFILL_83_DFFSR_125 gnd vdd FILL
XFILL_83_DFFSR_136 gnd vdd FILL
XFILL_83_DFFSR_147 gnd vdd FILL
XFILL_83_DFFSR_158 gnd vdd FILL
XFILL_83_DFFSR_169 gnd vdd FILL
XFILL_15_CLKBUF1_9 gnd vdd FILL
XFILL_3_DFFSR_206 gnd vdd FILL
XFILL_87_DFFSR_102 gnd vdd FILL
XFILL_0_NAND3X1_6 gnd vdd FILL
XFILL_3_DFFSR_217 gnd vdd FILL
XFILL_87_DFFSR_113 gnd vdd FILL
XFILL_87_DFFSR_124 gnd vdd FILL
XFILL_3_DFFSR_228 gnd vdd FILL
XFILL_87_DFFSR_135 gnd vdd FILL
XFILL_3_DFFSR_239 gnd vdd FILL
XFILL_87_DFFSR_146 gnd vdd FILL
XFILL_87_DFFSR_157 gnd vdd FILL
XFILL_23_DFFSR_19 gnd vdd FILL
XFILL_11_BUFX4_104 gnd vdd FILL
XFILL_14_BUFX4_40 gnd vdd FILL
XFILL_14_BUFX4_51 gnd vdd FILL
XFILL_87_DFFSR_168 gnd vdd FILL
XFILL_3_MUX2X1_180 gnd vdd FILL
XFILL_87_DFFSR_179 gnd vdd FILL
XFILL_19_CLKBUF1_8 gnd vdd FILL
XFILL_14_BUFX4_62 gnd vdd FILL
XFILL_3_MUX2X1_191 gnd vdd FILL
XFILL_7_DFFSR_205 gnd vdd FILL
XFILL_14_BUFX4_73 gnd vdd FILL
XFILL_4_NAND3X1_5 gnd vdd FILL
XFILL_14_BUFX4_84 gnd vdd FILL
XFILL_7_DFFSR_216 gnd vdd FILL
XDFFSR_230 INVX1_71/A CLKBUF1_26/Y DFFSR_25/R vdd MUX2X1_58/Y gnd vdd DFFSR
XFILL_14_BUFX4_95 gnd vdd FILL
XDFFSR_241 INVX1_55/A CLKBUF1_5/Y DFFSR_49/R vdd MUX2X1_42/Y gnd vdd DFFSR
XFILL_7_DFFSR_227 gnd vdd FILL
XFILL_7_DFFSR_238 gnd vdd FILL
XDFFSR_252 INVX1_49/A DFFSR_2/CLK BUFX4_50/Y vdd MUX2X1_36/Y gnd vdd DFFSR
XFILL_7_DFFSR_249 gnd vdd FILL
XDFFSR_263 INVX1_39/A DFFSR_9/CLK DFFSR_9/R vdd MUX2X1_26/Y gnd vdd DFFSR
XDFFSR_274 NOR2X1_6/A DFFSR_9/CLK DFFSR_9/R vdd DFFSR_274/D gnd vdd DFFSR
XFILL_63_DFFSR_18 gnd vdd FILL
XFILL_15_BUFX4_103 gnd vdd FILL
XFILL_63_DFFSR_29 gnd vdd FILL
XFILL_8_NAND3X1_4 gnd vdd FILL
XFILL_32_DFFSR_17 gnd vdd FILL
XFILL_32_DFFSR_28 gnd vdd FILL
XFILL_32_DFFSR_39 gnd vdd FILL
XFILL_57_5_1 gnd vdd FILL
XFILL_7_OAI22X1_18 gnd vdd FILL
XFILL_7_OAI22X1_29 gnd vdd FILL
XFILL_56_0_0 gnd vdd FILL
XFILL_72_DFFSR_190 gnd vdd FILL
XFILL_72_DFFSR_16 gnd vdd FILL
XFILL_23_DFFSR_203 gnd vdd FILL
XFILL_72_DFFSR_27 gnd vdd FILL
XFILL_72_DFFSR_38 gnd vdd FILL
XFILL_23_DFFSR_214 gnd vdd FILL
XFILL_72_DFFSR_49 gnd vdd FILL
XFILL_23_DFFSR_225 gnd vdd FILL
XFILL_23_DFFSR_236 gnd vdd FILL
XFILL_15_MUX2X1_6 gnd vdd FILL
XFILL_6_NAND3X1_50 gnd vdd FILL
XFILL_23_DFFSR_247 gnd vdd FILL
XFILL_6_NAND3X1_61 gnd vdd FILL
XFILL_23_DFFSR_258 gnd vdd FILL
XFILL_23_DFFSR_269 gnd vdd FILL
XFILL_6_NAND3X1_72 gnd vdd FILL
XFILL_27_DFFSR_202 gnd vdd FILL
XFILL_4_INVX1_209 gnd vdd FILL
XFILL_50_DFFSR_103 gnd vdd FILL
XFILL_6_NAND3X1_83 gnd vdd FILL
XFILL_6_NAND3X1_94 gnd vdd FILL
XFILL_50_DFFSR_114 gnd vdd FILL
XFILL_27_DFFSR_213 gnd vdd FILL
XFILL_50_DFFSR_125 gnd vdd FILL
XFILL_6_BUFX4_50 gnd vdd FILL
XFILL_27_DFFSR_224 gnd vdd FILL
XFILL_50_DFFSR_136 gnd vdd FILL
XFILL_27_DFFSR_235 gnd vdd FILL
XFILL_6_BUFX4_61 gnd vdd FILL
XFILL_8_AOI22X1_9 gnd vdd FILL
XFILL_41_DFFSR_15 gnd vdd FILL
XFILL_40_4_1 gnd vdd FILL
XFILL_6_BUFX4_72 gnd vdd FILL
XFILL_27_DFFSR_246 gnd vdd FILL
XFILL_50_DFFSR_147 gnd vdd FILL
XFILL_6_BUFX4_83 gnd vdd FILL
XFILL_50_DFFSR_158 gnd vdd FILL
XFILL_41_DFFSR_26 gnd vdd FILL
XFILL_41_DFFSR_37 gnd vdd FILL
XFILL_50_DFFSR_169 gnd vdd FILL
XFILL_27_DFFSR_257 gnd vdd FILL
XFILL_27_DFFSR_268 gnd vdd FILL
XFILL_41_DFFSR_48 gnd vdd FILL
XFILL_6_BUFX4_94 gnd vdd FILL
XFILL_41_DFFSR_59 gnd vdd FILL
XFILL_54_DFFSR_102 gnd vdd FILL
XFILL_18_CLKBUF1_16 gnd vdd FILL
XFILL_8_BUFX2_2 gnd vdd FILL
XFILL_54_DFFSR_113 gnd vdd FILL
XFILL_54_DFFSR_124 gnd vdd FILL
XFILL_18_CLKBUF1_27 gnd vdd FILL
XFILL_18_CLKBUF1_38 gnd vdd FILL
XFILL_54_DFFSR_135 gnd vdd FILL
XFILL_81_DFFSR_14 gnd vdd FILL
XFILL_54_DFFSR_146 gnd vdd FILL
XFILL_13_AOI21X1_13 gnd vdd FILL
XFILL_81_DFFSR_25 gnd vdd FILL
XFILL_54_DFFSR_157 gnd vdd FILL
XFILL_13_AOI21X1_24 gnd vdd FILL
XFILL_81_DFFSR_36 gnd vdd FILL
XFILL_54_DFFSR_168 gnd vdd FILL
XFILL_54_DFFSR_179 gnd vdd FILL
XFILL_13_AOI21X1_35 gnd vdd FILL
XFILL_81_DFFSR_47 gnd vdd FILL
XFILL_13_AOI21X1_46 gnd vdd FILL
XFILL_81_DFFSR_58 gnd vdd FILL
XFILL_10_DFFSR_14 gnd vdd FILL
XFILL_58_DFFSR_101 gnd vdd FILL
XFILL_13_AOI21X1_57 gnd vdd FILL
XFILL_81_DFFSR_69 gnd vdd FILL
XFILL_10_DFFSR_25 gnd vdd FILL
XFILL_13_AOI21X1_68 gnd vdd FILL
XFILL_58_DFFSR_112 gnd vdd FILL
XFILL_10_DFFSR_36 gnd vdd FILL
XFILL_13_AOI21X1_79 gnd vdd FILL
XFILL_58_DFFSR_123 gnd vdd FILL
XFILL_58_DFFSR_134 gnd vdd FILL
XFILL_10_DFFSR_47 gnd vdd FILL
XFILL_10_DFFSR_58 gnd vdd FILL
XFILL_67_DFFSR_1 gnd vdd FILL
XFILL_58_DFFSR_145 gnd vdd FILL
XFILL_10_DFFSR_69 gnd vdd FILL
XFILL_58_DFFSR_156 gnd vdd FILL
XFILL_8_NOR2X1_7 gnd vdd FILL
XFILL_58_DFFSR_167 gnd vdd FILL
XFILL_58_DFFSR_178 gnd vdd FILL
XFILL_50_DFFSR_13 gnd vdd FILL
XFILL_1_DFFSR_105 gnd vdd FILL
XFILL_58_DFFSR_189 gnd vdd FILL
XFILL_50_DFFSR_24 gnd vdd FILL
XFILL_1_DFFSR_116 gnd vdd FILL
XFILL_50_DFFSR_35 gnd vdd FILL
XFILL_1_DFFSR_127 gnd vdd FILL
XFILL_1_DFFSR_138 gnd vdd FILL
XFILL_50_DFFSR_46 gnd vdd FILL
XFILL_1_DFFSR_149 gnd vdd FILL
XFILL_50_DFFSR_57 gnd vdd FILL
XFILL_50_DFFSR_68 gnd vdd FILL
XFILL_50_DFFSR_79 gnd vdd FILL
XFILL_5_DFFSR_104 gnd vdd FILL
XFILL_48_5_1 gnd vdd FILL
XFILL_7_MUX2X1_5 gnd vdd FILL
XFILL_5_DFFSR_115 gnd vdd FILL
XFILL_5_DFFSR_126 gnd vdd FILL
XFILL_5_DFFSR_137 gnd vdd FILL
XFILL_47_0_0 gnd vdd FILL
XFILL_5_DFFSR_148 gnd vdd FILL
XFILL_25_CLKBUF1_40 gnd vdd FILL
XFILL_5_DFFSR_159 gnd vdd FILL
XFILL_51_DFFSR_7 gnd vdd FILL
XFILL_9_NAND3X1_107 gnd vdd FILL
XFILL_8_CLKBUF1_11 gnd vdd FILL
XFILL_9_NAND3X1_118 gnd vdd FILL
XFILL_9_DFFSR_103 gnd vdd FILL
XFILL_8_CLKBUF1_22 gnd vdd FILL
XFILL_9_NAND3X1_129 gnd vdd FILL
XFILL_9_DFFSR_114 gnd vdd FILL
XFILL_13_MUX2X1_12 gnd vdd FILL
XFILL_13_MUX2X1_23 gnd vdd FILL
XFILL_8_CLKBUF1_33 gnd vdd FILL
XFILL_9_DFFSR_125 gnd vdd FILL
XFILL_9_DFFSR_136 gnd vdd FILL
XFILL_13_MUX2X1_34 gnd vdd FILL
XFILL_16_MUX2X1_107 gnd vdd FILL
XFILL_16_MUX2X1_118 gnd vdd FILL
XFILL_13_MUX2X1_45 gnd vdd FILL
XFILL_9_DFFSR_147 gnd vdd FILL
XFILL_9_DFFSR_158 gnd vdd FILL
XFILL_16_MUX2X1_129 gnd vdd FILL
XFILL_3_AOI21X1_30 gnd vdd FILL
XFILL_13_MUX2X1_56 gnd vdd FILL
XFILL_3_AOI21X1_41 gnd vdd FILL
XFILL_9_DFFSR_169 gnd vdd FILL
XFILL_13_MUX2X1_67 gnd vdd FILL
XFILL_30_NOR3X1_8 gnd vdd FILL
XFILL_13_MUX2X1_78 gnd vdd FILL
XFILL_3_AOI21X1_52 gnd vdd FILL
XFILL_1_NOR3X1_16 gnd vdd FILL
XOAI21X1_11 INVX1_167/Y OAI21X1_2/B OAI21X1_11/C gnd NOR2X1_75/B vdd OAI21X1
XFILL_13_OAI22X1_10 gnd vdd FILL
XFILL_1_NOR3X1_27 gnd vdd FILL
XFILL_13_MUX2X1_89 gnd vdd FILL
XOAI21X1_22 INVX1_148/Y OAI21X1_4/B OAI21X1_22/C gnd NOR2X1_93/A vdd OAI21X1
XFILL_3_AOI21X1_63 gnd vdd FILL
XFILL_13_OAI22X1_21 gnd vdd FILL
XFILL_3_AOI21X1_74 gnd vdd FILL
XFILL_1_NOR3X1_38 gnd vdd FILL
XFILL_13_OAI22X1_32 gnd vdd FILL
XFILL_17_MUX2X1_11 gnd vdd FILL
XFILL_17_MUX2X1_22 gnd vdd FILL
XFILL_1_NOR3X1_49 gnd vdd FILL
XOAI21X1_33 NOR2X1_24/A OAI21X1_46/B AOI22X1_3/A gnd OAI21X1_33/Y vdd OAI21X1
XFILL_31_4_1 gnd vdd FILL
XFILL_13_OAI22X1_43 gnd vdd FILL
XOAI21X1_44 INVX2_3/Y NOR2X1_24/A NOR2X1_13/B gnd OAI21X1_46/C vdd OAI21X1
XFILL_17_MUX2X1_33 gnd vdd FILL
XFILL_17_MUX2X1_44 gnd vdd FILL
XFILL_17_MUX2X1_55 gnd vdd FILL
XFILL_2_DFFSR_13 gnd vdd FILL
XFILL_17_MUX2X1_66 gnd vdd FILL
XFILL_6_NOR2X1_140 gnd vdd FILL
XFILL_17_MUX2X1_77 gnd vdd FILL
XFILL_2_DFFSR_24 gnd vdd FILL
XFILL_17_MUX2X1_88 gnd vdd FILL
XFILL_2_DFFSR_35 gnd vdd FILL
XFILL_5_NOR3X1_15 gnd vdd FILL
XFILL_6_NOR2X1_151 gnd vdd FILL
XFILL_5_NOR3X1_26 gnd vdd FILL
XFILL_6_NOR2X1_162 gnd vdd FILL
XFILL_2_DFFSR_46 gnd vdd FILL
XFILL_13_NAND3X1_120 gnd vdd FILL
XFILL_17_MUX2X1_99 gnd vdd FILL
XFILL_13_NAND3X1_131 gnd vdd FILL
XFILL_6_NOR2X1_173 gnd vdd FILL
XFILL_5_NOR3X1_37 gnd vdd FILL
XFILL_21_DFFSR_102 gnd vdd FILL
XFILL_2_DFFSR_57 gnd vdd FILL
XFILL_6_NOR2X1_184 gnd vdd FILL
XFILL_5_NOR3X1_48 gnd vdd FILL
XFILL_2_DFFSR_68 gnd vdd FILL
XFILL_6_NOR2X1_195 gnd vdd FILL
XFILL_21_DFFSR_113 gnd vdd FILL
XFILL_21_DFFSR_124 gnd vdd FILL
XFILL_2_DFFSR_79 gnd vdd FILL
XFILL_21_DFFSR_135 gnd vdd FILL
XFILL_21_DFFSR_146 gnd vdd FILL
XFILL_10_NOR2X1_201 gnd vdd FILL
XFILL_21_DFFSR_157 gnd vdd FILL
XFILL_9_NOR3X1_14 gnd vdd FILL
XFILL_21_DFFSR_168 gnd vdd FILL
XFILL_21_DFFSR_179 gnd vdd FILL
XFILL_9_NOR3X1_25 gnd vdd FILL
XFILL_2_INVX1_108 gnd vdd FILL
XFILL_9_NOR3X1_36 gnd vdd FILL
XFILL_25_DFFSR_101 gnd vdd FILL
XFILL_9_NOR3X1_47 gnd vdd FILL
XFILL_2_INVX1_119 gnd vdd FILL
XFILL_25_DFFSR_112 gnd vdd FILL
XFILL_25_DFFSR_123 gnd vdd FILL
XFILL_25_DFFSR_134 gnd vdd FILL
XFILL_23_MUX2X1_120 gnd vdd FILL
XFILL_25_DFFSR_145 gnd vdd FILL
XFILL_23_MUX2X1_131 gnd vdd FILL
XFILL_25_DFFSR_156 gnd vdd FILL
XFILL_4_NAND3X1_103 gnd vdd FILL
XFILL_4_NAND3X1_114 gnd vdd FILL
XFILL_25_DFFSR_167 gnd vdd FILL
XFILL_23_MUX2X1_142 gnd vdd FILL
XFILL_25_DFFSR_178 gnd vdd FILL
XFILL_23_MUX2X1_153 gnd vdd FILL
XFILL_4_NAND3X1_125 gnd vdd FILL
XFILL_6_INVX1_107 gnd vdd FILL
XFILL_6_MUX2X1_102 gnd vdd FILL
XFILL_23_MUX2X1_164 gnd vdd FILL
XFILL_23_MUX2X1_175 gnd vdd FILL
XFILL_6_INVX1_118 gnd vdd FILL
XFILL_29_DFFSR_100 gnd vdd FILL
XFILL_25_DFFSR_189 gnd vdd FILL
XFILL_6_MUX2X1_113 gnd vdd FILL
XFILL_6_INVX1_129 gnd vdd FILL
XFILL_23_MUX2X1_186 gnd vdd FILL
XFILL_29_DFFSR_111 gnd vdd FILL
XFILL_6_MUX2X1_124 gnd vdd FILL
XFILL_29_DFFSR_122 gnd vdd FILL
XFILL_29_DFFSR_133 gnd vdd FILL
XFILL_6_MUX2X1_135 gnd vdd FILL
XFILL_6_MUX2X1_146 gnd vdd FILL
XFILL_29_DFFSR_144 gnd vdd FILL
XFILL_6_MUX2X1_157 gnd vdd FILL
XFILL_29_DFFSR_155 gnd vdd FILL
XFILL_39_5_1 gnd vdd FILL
XFILL_6_MUX2X1_168 gnd vdd FILL
XFILL_29_DFFSR_166 gnd vdd FILL
XFILL_19_DFFSR_80 gnd vdd FILL
XFILL_29_DFFSR_177 gnd vdd FILL
XFILL_6_MUX2X1_179 gnd vdd FILL
XFILL_21_NOR3X1_13 gnd vdd FILL
XFILL_38_0_0 gnd vdd FILL
XFILL_19_DFFSR_91 gnd vdd FILL
XFILL_29_DFFSR_188 gnd vdd FILL
XFILL_21_NOR3X1_24 gnd vdd FILL
XFILL_21_NOR3X1_35 gnd vdd FILL
XFILL_29_DFFSR_199 gnd vdd FILL
XFILL_21_NOR3X1_46 gnd vdd FILL
XFILL_71_DFFSR_202 gnd vdd FILL
XFILL_71_DFFSR_213 gnd vdd FILL
XFILL_7_OAI21X1_40 gnd vdd FILL
XFILL_71_DFFSR_224 gnd vdd FILL
XFILL_71_DFFSR_235 gnd vdd FILL
XFILL_71_DFFSR_246 gnd vdd FILL
XFILL_25_NOR3X1_12 gnd vdd FILL
XFILL_59_DFFSR_90 gnd vdd FILL
XFILL_71_DFFSR_257 gnd vdd FILL
XFILL_71_DFFSR_268 gnd vdd FILL
XFILL_25_NOR3X1_23 gnd vdd FILL
XFILL_25_NOR3X1_34 gnd vdd FILL
XFILL_75_DFFSR_201 gnd vdd FILL
XFILL_25_NOR3X1_45 gnd vdd FILL
XFILL_75_DFFSR_212 gnd vdd FILL
XFILL_75_DFFSR_223 gnd vdd FILL
XFILL_75_DFFSR_234 gnd vdd FILL
XFILL_22_4_1 gnd vdd FILL
XFILL_75_DFFSR_245 gnd vdd FILL
XFILL_29_NOR3X1_11 gnd vdd FILL
XFILL_75_DFFSR_256 gnd vdd FILL
XFILL_29_NOR3X1_22 gnd vdd FILL
XFILL_75_DFFSR_267 gnd vdd FILL
XFILL_29_NOR3X1_33 gnd vdd FILL
XFILL_30_CLKBUF1_8 gnd vdd FILL
XFILL_79_DFFSR_200 gnd vdd FILL
XFILL_29_NOR3X1_44 gnd vdd FILL
XFILL_79_DFFSR_211 gnd vdd FILL
XFILL_79_DFFSR_222 gnd vdd FILL
XFILL_79_DFFSR_233 gnd vdd FILL
XFILL_79_DFFSR_244 gnd vdd FILL
XFILL_79_DFFSR_255 gnd vdd FILL
XFILL_34_CLKBUF1_7 gnd vdd FILL
XFILL_79_DFFSR_266 gnd vdd FILL
XFILL_9_NAND3X1_16 gnd vdd FILL
XFILL_9_NAND3X1_27 gnd vdd FILL
XFILL_9_NAND3X1_38 gnd vdd FILL
XFILL_9_NAND3X1_49 gnd vdd FILL
XFILL_15_BUFX4_18 gnd vdd FILL
XFILL_15_BUFX4_29 gnd vdd FILL
XFILL_0_NOR3X1_4 gnd vdd FILL
XFILL_5_5_1 gnd vdd FILL
XFILL_29_0_0 gnd vdd FILL
XFILL_4_0_0 gnd vdd FILL
XFILL_2_NAND2X1_18 gnd vdd FILL
XFILL_33_DFFSR_4 gnd vdd FILL
XFILL_2_NAND2X1_29 gnd vdd FILL
XFILL_0_OAI21X1_3 gnd vdd FILL
XFILL_12_MUX2X1_160 gnd vdd FILL
XFILL_12_MUX2X1_171 gnd vdd FILL
XFILL_12_MUX2X1_182 gnd vdd FILL
XFILL_13_4_1 gnd vdd FILL
XFILL_12_MUX2X1_193 gnd vdd FILL
XFILL_42_DFFSR_201 gnd vdd FILL
XFILL_42_DFFSR_212 gnd vdd FILL
XFILL_4_OAI21X1_2 gnd vdd FILL
XFILL_42_DFFSR_223 gnd vdd FILL
XFILL_42_DFFSR_234 gnd vdd FILL
XFILL_42_DFFSR_245 gnd vdd FILL
XFILL_1_NOR2X1_60 gnd vdd FILL
XFILL_1_NOR2X1_71 gnd vdd FILL
XFILL_42_DFFSR_256 gnd vdd FILL
XFILL_42_DFFSR_267 gnd vdd FILL
XFILL_1_NOR2X1_82 gnd vdd FILL
XFILL_1_NOR2X1_93 gnd vdd FILL
XFILL_46_DFFSR_200 gnd vdd FILL
XFILL_28_CLKBUF1_17 gnd vdd FILL
XFILL_28_CLKBUF1_28 gnd vdd FILL
XFILL_46_DFFSR_211 gnd vdd FILL
XFILL_8_OAI21X1_1 gnd vdd FILL
XFILL_46_DFFSR_222 gnd vdd FILL
XFILL_28_CLKBUF1_39 gnd vdd FILL
XFILL_46_DFFSR_233 gnd vdd FILL
XFILL_7_BUFX4_17 gnd vdd FILL
XFILL_55_DFFSR_8 gnd vdd FILL
XFILL_46_DFFSR_244 gnd vdd FILL
XFILL_7_BUFX4_28 gnd vdd FILL
XFILL_46_DFFSR_255 gnd vdd FILL
XFILL_7_BUFX4_39 gnd vdd FILL
XFILL_5_NOR2X1_70 gnd vdd FILL
XFILL_5_NOR2X1_81 gnd vdd FILL
XFILL_46_DFFSR_266 gnd vdd FILL
XFILL_5_NOR2X1_92 gnd vdd FILL
XFILL_73_DFFSR_100 gnd vdd FILL
XFILL_73_DFFSR_111 gnd vdd FILL
XFILL_73_DFFSR_122 gnd vdd FILL
XFILL_6_AOI21X1_18 gnd vdd FILL
XFILL_73_DFFSR_133 gnd vdd FILL
XFILL_6_AOI21X1_29 gnd vdd FILL
XFILL_73_DFFSR_144 gnd vdd FILL
XFILL_73_DFFSR_155 gnd vdd FILL
XFILL_73_DFFSR_166 gnd vdd FILL
XFILL_73_DFFSR_177 gnd vdd FILL
XFILL_9_NOR2X1_80 gnd vdd FILL
XFILL_73_DFFSR_188 gnd vdd FILL
XFILL_9_NOR2X1_91 gnd vdd FILL
XFILL_6_4 gnd vdd FILL
XFILL_77_DFFSR_110 gnd vdd FILL
XFILL_73_DFFSR_199 gnd vdd FILL
XFILL_9_NOR2X1_106 gnd vdd FILL
XFILL_77_DFFSR_121 gnd vdd FILL
XFILL_77_DFFSR_132 gnd vdd FILL
XFILL_9_NOR2X1_117 gnd vdd FILL
XFILL_77_DFFSR_143 gnd vdd FILL
XFILL_9_NOR2X1_128 gnd vdd FILL
XFILL_9_NOR2X1_139 gnd vdd FILL
XFILL_77_DFFSR_154 gnd vdd FILL
XFILL_77_DFFSR_165 gnd vdd FILL
XFILL_15_NAND3X1_30 gnd vdd FILL
XFILL_15_NAND3X1_41 gnd vdd FILL
XFILL_77_DFFSR_176 gnd vdd FILL
XFILL_77_DFFSR_187 gnd vdd FILL
XFILL_15_NAND3X1_52 gnd vdd FILL
XFILL_15_NAND3X1_63 gnd vdd FILL
XFILL_77_DFFSR_198 gnd vdd FILL
XFILL_15_NAND3X1_74 gnd vdd FILL
XFILL_14_AND2X2_5 gnd vdd FILL
XFILL_35_CLKBUF1_30 gnd vdd FILL
XFILL_15_NAND3X1_85 gnd vdd FILL
XFILL_35_CLKBUF1_41 gnd vdd FILL
XFILL_15_NAND3X1_96 gnd vdd FILL
XFILL_63_3_1 gnd vdd FILL
XFILL_1_NAND2X1_4 gnd vdd FILL
XFILL_11_BUFX4_11 gnd vdd FILL
XFILL_11_BUFX4_22 gnd vdd FILL
XFILL_11_BUFX4_33 gnd vdd FILL
XFILL_11_BUFX4_44 gnd vdd FILL
XFILL_5_NAND2X1_3 gnd vdd FILL
XFILL_11_BUFX4_55 gnd vdd FILL
XFILL_11_BUFX4_66 gnd vdd FILL
XFILL_11_BUFX4_77 gnd vdd FILL
XFILL_11_BUFX4_88 gnd vdd FILL
XFILL_11_BUFX4_99 gnd vdd FILL
XFILL_6_OAI22X1_15 gnd vdd FILL
XFILL_6_OAI22X1_26 gnd vdd FILL
XFILL_6_OAI22X1_37 gnd vdd FILL
XFILL_14_NAND3X1_110 gnd vdd FILL
XFILL_14_NAND3X1_121 gnd vdd FILL
XDFFSR_14 INVX1_33/A DFFSR_7/CLK DFFSR_26/R vdd DFFSR_14/D gnd vdd DFFSR
XFILL_6_OAI22X1_48 gnd vdd FILL
XFILL_14_NAND3X1_132 gnd vdd FILL
XDFFSR_25 DFFSR_25/Q DFFSR_87/CLK DFFSR_25/R vdd DFFSR_25/D gnd vdd DFFSR
XFILL_9_NAND2X1_2 gnd vdd FILL
XFILL_13_DFFSR_200 gnd vdd FILL
XDFFSR_36 DFFSR_36/Q DFFSR_47/CLK DFFSR_79/R vdd DFFSR_36/D gnd vdd DFFSR
XFILL_13_DFFSR_211 gnd vdd FILL
XDFFSR_47 INVX1_14/A DFFSR_47/CLK DFFSR_79/R vdd DFFSR_47/D gnd vdd DFFSR
XFILL_13_DFFSR_222 gnd vdd FILL
XDFFSR_58 INVX1_6/A DFFSR_58/CLK DFFSR_58/R vdd DFFSR_58/D gnd vdd DFFSR
XFILL_13_DFFSR_233 gnd vdd FILL
XDFFSR_69 DFFSR_69/Q DFFSR_73/CLK DFFSR_69/R vdd DFFSR_69/D gnd vdd DFFSR
XFILL_13_DFFSR_244 gnd vdd FILL
XFILL_13_DFFSR_255 gnd vdd FILL
XFILL_13_DFFSR_266 gnd vdd FILL
XFILL_5_NAND3X1_80 gnd vdd FILL
XFILL_40_DFFSR_100 gnd vdd FILL
XFILL_5_NAND3X1_91 gnd vdd FILL
XFILL_17_DFFSR_210 gnd vdd FILL
XFILL_40_DFFSR_111 gnd vdd FILL
XFILL_9_NAND2X1_60 gnd vdd FILL
XFILL_3_NOR2X1_206 gnd vdd FILL
XFILL_40_DFFSR_122 gnd vdd FILL
XFILL_17_DFFSR_221 gnd vdd FILL
XFILL_1_AOI21X1_9 gnd vdd FILL
XFILL_40_DFFSR_133 gnd vdd FILL
XFILL_17_DFFSR_232 gnd vdd FILL
XFILL_9_NAND2X1_71 gnd vdd FILL
XFILL_5_INVX1_12 gnd vdd FILL
XFILL_17_DFFSR_243 gnd vdd FILL
XFILL_40_DFFSR_144 gnd vdd FILL
XFILL_5_INVX1_23 gnd vdd FILL
XFILL_9_NAND2X1_82 gnd vdd FILL
XCLKBUF1_12 BUFX4_10/Y gnd DFFSR_55/CLK vdd CLKBUF1
XFILL_5_INVX1_34 gnd vdd FILL
XFILL_40_DFFSR_155 gnd vdd FILL
XFILL_17_DFFSR_254 gnd vdd FILL
XFILL_9_NAND2X1_93 gnd vdd FILL
XFILL_5_NAND3X1_104 gnd vdd FILL
XCLKBUF1_23 BUFX4_73/Y gnd DFFSR_73/CLK vdd CLKBUF1
XFILL_5_NAND3X1_115 gnd vdd FILL
XFILL_5_INVX1_45 gnd vdd FILL
XFILL_40_DFFSR_166 gnd vdd FILL
XFILL_40_DFFSR_177 gnd vdd FILL
XFILL_6_AND2X2_4 gnd vdd FILL
XCLKBUF1_34 BUFX4_73/Y gnd CLKBUF1_34/Y vdd CLKBUF1
XFILL_5_NAND3X1_126 gnd vdd FILL
XFILL_17_DFFSR_265 gnd vdd FILL
XFILL_5_INVX1_56 gnd vdd FILL
XFILL_5_INVX1_67 gnd vdd FILL
XFILL_40_DFFSR_188 gnd vdd FILL
XFILL_5_INVX1_78 gnd vdd FILL
XFILL_44_DFFSR_110 gnd vdd FILL
XFILL_40_DFFSR_199 gnd vdd FILL
XFILL_17_CLKBUF1_13 gnd vdd FILL
XFILL_5_INVX1_89 gnd vdd FILL
XFILL_17_CLKBUF1_24 gnd vdd FILL
XFILL_44_DFFSR_121 gnd vdd FILL
XFILL_44_DFFSR_132 gnd vdd FILL
XFILL_17_CLKBUF1_35 gnd vdd FILL
XFILL_5_AOI21X1_8 gnd vdd FILL
XFILL_44_DFFSR_143 gnd vdd FILL
XFILL_12_AOI21X1_10 gnd vdd FILL
XFILL_44_DFFSR_154 gnd vdd FILL
XFILL_12_AOI21X1_21 gnd vdd FILL
XFILL_12_AOI21X1_32 gnd vdd FILL
XFILL_44_DFFSR_165 gnd vdd FILL
XFILL_44_DFFSR_176 gnd vdd FILL
XFILL_2_DFFSR_3 gnd vdd FILL
XFILL_12_AOI21X1_43 gnd vdd FILL
XFILL_44_DFFSR_187 gnd vdd FILL
XFILL_12_AOI21X1_54 gnd vdd FILL
XFILL_54_3_1 gnd vdd FILL
XFILL_44_DFFSR_198 gnd vdd FILL
XFILL_15_DFFSR_1 gnd vdd FILL
XFILL_12_AOI21X1_65 gnd vdd FILL
XFILL_3_BUFX4_10 gnd vdd FILL
XFILL_48_DFFSR_120 gnd vdd FILL
XFILL_12_AOI21X1_76 gnd vdd FILL
XFILL_48_DFFSR_131 gnd vdd FILL
XFILL_9_AOI21X1_7 gnd vdd FILL
XFILL_3_BUFX4_21 gnd vdd FILL
XFILL_72_DFFSR_2 gnd vdd FILL
XFILL_48_DFFSR_142 gnd vdd FILL
XFILL_3_BUFX4_32 gnd vdd FILL
XFILL_48_DFFSR_153 gnd vdd FILL
XFILL_3_BUFX4_43 gnd vdd FILL
XFILL_10_AOI22X1_5 gnd vdd FILL
XFILL_3_BUFX4_54 gnd vdd FILL
XFILL_48_DFFSR_164 gnd vdd FILL
XFILL_48_DFFSR_175 gnd vdd FILL
XFILL_3_BUFX4_65 gnd vdd FILL
XFILL_3_BUFX4_76 gnd vdd FILL
XFILL_48_DFFSR_186 gnd vdd FILL
XFILL_48_DFFSR_197 gnd vdd FILL
XFILL_3_BUFX4_87 gnd vdd FILL
XFILL_3_BUFX4_98 gnd vdd FILL
XFILL_10_BUFX2_7 gnd vdd FILL
XFILL_14_AOI22X1_4 gnd vdd FILL
XFILL_21_MUX2X1_8 gnd vdd FILL
XFILL_18_AOI22X1_3 gnd vdd FILL
XFILL_0_NAND3X1_100 gnd vdd FILL
XFILL_0_NAND3X1_111 gnd vdd FILL
XFILL_0_NAND3X1_122 gnd vdd FILL
XFILL_37_DFFSR_5 gnd vdd FILL
XINVX1_108 INVX1_108/A gnd MUX2X1_95/A vdd INVX1
XINVX1_119 NOR2X1_44/B gnd NAND3X1_2/C vdd INVX1
XFILL_7_CLKBUF1_30 gnd vdd FILL
XFILL_29_DFFSR_12 gnd vdd FILL
XFILL_7_CLKBUF1_41 gnd vdd FILL
XFILL_29_DFFSR_23 gnd vdd FILL
XFILL_15_MUX2X1_104 gnd vdd FILL
XFILL_29_DFFSR_34 gnd vdd FILL
XFILL_15_MUX2X1_115 gnd vdd FILL
XFILL_29_DFFSR_45 gnd vdd FILL
XFILL_15_MUX2X1_126 gnd vdd FILL
XFILL_29_DFFSR_56 gnd vdd FILL
XFILL_15_MUX2X1_137 gnd vdd FILL
XFILL_29_DFFSR_67 gnd vdd FILL
XFILL_29_DFFSR_78 gnd vdd FILL
XFILL_15_MUX2X1_148 gnd vdd FILL
XFILL_2_AOI21X1_60 gnd vdd FILL
XFILL_29_DFFSR_89 gnd vdd FILL
XFILL_15_MUX2X1_159 gnd vdd FILL
XFILL_2_AOI21X1_71 gnd vdd FILL
XFILL_69_DFFSR_11 gnd vdd FILL
XFILL_12_OAI22X1_40 gnd vdd FILL
XFILL_69_DFFSR_22 gnd vdd FILL
XFILL_12_OAI22X1_51 gnd vdd FILL
XFILL_69_DFFSR_33 gnd vdd FILL
XFILL_69_DFFSR_44 gnd vdd FILL
XFILL_4_MUX2X1_9 gnd vdd FILL
XFILL_69_DFFSR_55 gnd vdd FILL
XFILL_69_DFFSR_66 gnd vdd FILL
XFILL_69_DFFSR_77 gnd vdd FILL
XFILL_69_DFFSR_88 gnd vdd FILL
XFILL_69_DFFSR_99 gnd vdd FILL
XFILL_5_NOR2X1_170 gnd vdd FILL
XFILL_5_NOR2X1_181 gnd vdd FILL
XFILL_11_DFFSR_110 gnd vdd FILL
XFILL_5_NOR2X1_192 gnd vdd FILL
XFILL_11_DFFSR_121 gnd vdd FILL
XFILL_11_DFFSR_132 gnd vdd FILL
XFILL_59_DFFSR_9 gnd vdd FILL
XFILL_38_DFFSR_10 gnd vdd FILL
XFILL_11_DFFSR_143 gnd vdd FILL
XFILL_11_DFFSR_154 gnd vdd FILL
XFILL_38_DFFSR_21 gnd vdd FILL
XFILL_45_3_1 gnd vdd FILL
XFILL_11_DFFSR_165 gnd vdd FILL
XFILL_38_DFFSR_32 gnd vdd FILL
XFILL_38_DFFSR_43 gnd vdd FILL
XFILL_11_DFFSR_176 gnd vdd FILL
XFILL_0_CLKBUF1_8 gnd vdd FILL
XFILL_38_DFFSR_54 gnd vdd FILL
XFILL_38_DFFSR_65 gnd vdd FILL
XFILL_11_DFFSR_187 gnd vdd FILL
XFILL_11_DFFSR_198 gnd vdd FILL
XFILL_38_DFFSR_76 gnd vdd FILL
XFILL_15_DFFSR_120 gnd vdd FILL
XFILL_15_DFFSR_131 gnd vdd FILL
XFILL_38_DFFSR_87 gnd vdd FILL
XFILL_38_DFFSR_98 gnd vdd FILL
XFILL_15_DFFSR_142 gnd vdd FILL
XFILL_78_DFFSR_20 gnd vdd FILL
XFILL_15_DFFSR_153 gnd vdd FILL
XFILL_27_9 gnd vdd FILL
XFILL_78_DFFSR_31 gnd vdd FILL
XFILL_15_DFFSR_164 gnd vdd FILL
XFILL_4_CLKBUF1_7 gnd vdd FILL
XFILL_15_DFFSR_175 gnd vdd FILL
XFILL_22_MUX2X1_150 gnd vdd FILL
XFILL_78_DFFSR_42 gnd vdd FILL
XFILL_22_MUX2X1_161 gnd vdd FILL
XFILL_15_DFFSR_186 gnd vdd FILL
XFILL_78_DFFSR_53 gnd vdd FILL
XFILL_5_MUX2X1_110 gnd vdd FILL
XFILL_22_MUX2X1_172 gnd vdd FILL
XFILL_78_DFFSR_64 gnd vdd FILL
XFILL_15_DFFSR_197 gnd vdd FILL
XFILL_78_DFFSR_75 gnd vdd FILL
XFILL_22_MUX2X1_183 gnd vdd FILL
XFILL_5_MUX2X1_121 gnd vdd FILL
XFILL_22_MUX2X1_194 gnd vdd FILL
XFILL_19_DFFSR_130 gnd vdd FILL
XFILL_78_DFFSR_86 gnd vdd FILL
XFILL_5_MUX2X1_132 gnd vdd FILL
XFILL_5_MUX2X1_143 gnd vdd FILL
XFILL_19_DFFSR_141 gnd vdd FILL
XFILL_78_DFFSR_97 gnd vdd FILL
XFILL_5_MUX2X1_154 gnd vdd FILL
XFILL_19_DFFSR_152 gnd vdd FILL
XFILL_5_MUX2X1_165 gnd vdd FILL
XFILL_0_BUFX4_102 gnd vdd FILL
XFILL_1_INVX1_60 gnd vdd FILL
XFILL_19_DFFSR_163 gnd vdd FILL
XFILL_19_DFFSR_174 gnd vdd FILL
XFILL_11_NOR3X1_10 gnd vdd FILL
XFILL_5_MUX2X1_176 gnd vdd FILL
XFILL_8_CLKBUF1_6 gnd vdd FILL
XFILL_5_MUX2X1_187 gnd vdd FILL
XFILL_1_INVX1_71 gnd vdd FILL
XFILL_19_DFFSR_185 gnd vdd FILL
XFILL_1_INVX1_82 gnd vdd FILL
XFILL_11_NOR3X1_21 gnd vdd FILL
XFILL_19_DFFSR_196 gnd vdd FILL
XFILL_1_INVX1_93 gnd vdd FILL
XFILL_47_DFFSR_30 gnd vdd FILL
XFILL_11_NOR3X1_32 gnd vdd FILL
XFILL_11_NOR3X1_43 gnd vdd FILL
XFILL_18_NOR3X1_5 gnd vdd FILL
XFILL_47_DFFSR_41 gnd vdd FILL
XFILL_61_DFFSR_210 gnd vdd FILL
XFILL_47_DFFSR_52 gnd vdd FILL
XFILL_47_DFFSR_63 gnd vdd FILL
XFILL_61_DFFSR_221 gnd vdd FILL
XFILL_4_BUFX4_101 gnd vdd FILL
XFILL_47_DFFSR_74 gnd vdd FILL
XFILL_61_DFFSR_232 gnd vdd FILL
XFILL_61_DFFSR_243 gnd vdd FILL
XFILL_47_DFFSR_85 gnd vdd FILL
XFILL_61_DFFSR_254 gnd vdd FILL
XFILL_47_DFFSR_96 gnd vdd FILL
XFILL_15_NOR3X1_20 gnd vdd FILL
XFILL_61_DFFSR_265 gnd vdd FILL
XFILL_15_NOR3X1_31 gnd vdd FILL
XFILL_87_DFFSR_40 gnd vdd FILL
XFILL_15_NOR3X1_42 gnd vdd FILL
XFILL_87_DFFSR_51 gnd vdd FILL
XFILL_87_DFFSR_62 gnd vdd FILL
XFILL_65_DFFSR_220 gnd vdd FILL
XFILL_8_BUFX4_100 gnd vdd FILL
XFILL_87_DFFSR_73 gnd vdd FILL
XFILL_65_DFFSR_231 gnd vdd FILL
XFILL_87_DFFSR_84 gnd vdd FILL
XFILL_16_DFFSR_40 gnd vdd FILL
XFILL_65_DFFSR_242 gnd vdd FILL
XFILL_87_DFFSR_95 gnd vdd FILL
XFILL_4_1 gnd vdd FILL
XFILL_65_DFFSR_253 gnd vdd FILL
XFILL_16_DFFSR_51 gnd vdd FILL
XFILL_65_DFFSR_264 gnd vdd FILL
XFILL_16_DFFSR_62 gnd vdd FILL
XFILL_20_CLKBUF1_5 gnd vdd FILL
XFILL_65_DFFSR_275 gnd vdd FILL
XFILL_16_DFFSR_73 gnd vdd FILL
XFILL_19_NOR3X1_30 gnd vdd FILL
XFILL_16_DFFSR_84 gnd vdd FILL
XFILL_19_NOR3X1_41 gnd vdd FILL
XFILL_16_DFFSR_95 gnd vdd FILL
XFILL_19_NOR3X1_52 gnd vdd FILL
XFILL_60_3 gnd vdd FILL
XFILL_69_DFFSR_230 gnd vdd FILL
XFILL_27_NOR3X1_3 gnd vdd FILL
XFILL_69_DFFSR_241 gnd vdd FILL
XFILL_53_2 gnd vdd FILL
XFILL_69_DFFSR_252 gnd vdd FILL
XFILL_56_DFFSR_50 gnd vdd FILL
XFILL_69_DFFSR_263 gnd vdd FILL
XFILL_24_CLKBUF1_4 gnd vdd FILL
XFILL_56_DFFSR_61 gnd vdd FILL
XFILL_69_DFFSR_274 gnd vdd FILL
XFILL_56_DFFSR_72 gnd vdd FILL
XFILL_56_DFFSR_83 gnd vdd FILL
XFILL_46_1 gnd vdd FILL
XFILL_36_3_1 gnd vdd FILL
XFILL_56_DFFSR_94 gnd vdd FILL
XFILL_2_NOR2X1_14 gnd vdd FILL
XFILL_2_NOR2X1_25 gnd vdd FILL
XFILL_8_NAND3X1_13 gnd vdd FILL
XFILL_2_NOR2X1_36 gnd vdd FILL
XFILL_8_NAND3X1_24 gnd vdd FILL
XFILL_2_NOR2X1_47 gnd vdd FILL
XFILL_8_NAND3X1_35 gnd vdd FILL
XFILL_1_NOR2X1_4 gnd vdd FILL
XFILL_2_NOR2X1_58 gnd vdd FILL
XFILL_8_NAND3X1_46 gnd vdd FILL
XFILL_8_NAND3X1_57 gnd vdd FILL
XFILL_2_NOR2X1_69 gnd vdd FILL
XFILL_28_CLKBUF1_3 gnd vdd FILL
XFILL_8_NAND3X1_68 gnd vdd FILL
XFILL_8_NAND3X1_79 gnd vdd FILL
XFILL_6_NOR2X1_13 gnd vdd FILL
XFILL_47_DFFSR_209 gnd vdd FILL
XFILL_25_DFFSR_60 gnd vdd FILL
XFILL_6_NOR2X1_24 gnd vdd FILL
XFILL_6_NOR2X1_35 gnd vdd FILL
XFILL_25_DFFSR_71 gnd vdd FILL
XFILL_6_NOR2X1_46 gnd vdd FILL
XFILL_25_DFFSR_82 gnd vdd FILL
XFILL_10_OAI22X1_8 gnd vdd FILL
XFILL_25_DFFSR_93 gnd vdd FILL
XFILL_6_NOR2X1_57 gnd vdd FILL
XFILL_6_NOR2X1_68 gnd vdd FILL
XFILL_6_NOR2X1_79 gnd vdd FILL
XFILL_20_7_2 gnd vdd FILL
XFILL_0_MUX2X1_2 gnd vdd FILL
XFILL_74_DFFSR_109 gnd vdd FILL
XFILL_65_DFFSR_70 gnd vdd FILL
XFILL_65_DFFSR_81 gnd vdd FILL
XFILL_65_DFFSR_92 gnd vdd FILL
XFILL_14_OAI22X1_7 gnd vdd FILL
XFILL_15_NAND3X1_100 gnd vdd FILL
XFILL_15_NAND3X1_111 gnd vdd FILL
XFILL_1_NAND2X1_15 gnd vdd FILL
XFILL_6_DFFSR_4 gnd vdd FILL
XFILL_1_NAND2X1_26 gnd vdd FILL
XFILL_1_NAND2X1_37 gnd vdd FILL
XFILL_15_NAND3X1_122 gnd vdd FILL
XFILL_1_NAND2X1_48 gnd vdd FILL
XFILL_19_DFFSR_2 gnd vdd FILL
XFILL_78_DFFSR_108 gnd vdd FILL
XFILL_1_NAND2X1_59 gnd vdd FILL
XFILL_76_DFFSR_3 gnd vdd FILL
XFILL_78_DFFSR_119 gnd vdd FILL
XFILL_8_DFFSR_50 gnd vdd FILL
XFILL_8_DFFSR_61 gnd vdd FILL
XFILL_18_OAI22X1_6 gnd vdd FILL
XFILL_8_DFFSR_72 gnd vdd FILL
XFILL_8_DFFSR_83 gnd vdd FILL
XFILL_8_DFFSR_94 gnd vdd FILL
XFILL_34_DFFSR_80 gnd vdd FILL
XFILL_11_MUX2X1_190 gnd vdd FILL
XFILL_34_DFFSR_91 gnd vdd FILL
XFILL_32_DFFSR_220 gnd vdd FILL
XFILL_32_DFFSR_231 gnd vdd FILL
XFILL_32_DFFSR_242 gnd vdd FILL
XFILL_32_DFFSR_253 gnd vdd FILL
XFILL_6_NAND3X1_105 gnd vdd FILL
XFILL_6_NAND3X1_116 gnd vdd FILL
XFILL_32_DFFSR_264 gnd vdd FILL
XFILL_6_NAND3X1_127 gnd vdd FILL
XFILL_32_DFFSR_275 gnd vdd FILL
XFILL_74_DFFSR_90 gnd vdd FILL
XFILL_27_CLKBUF1_14 gnd vdd FILL
XFILL_27_CLKBUF1_25 gnd vdd FILL
XFILL_27_CLKBUF1_36 gnd vdd FILL
XFILL_60_DFFSR_9 gnd vdd FILL
XFILL_36_DFFSR_230 gnd vdd FILL
XFILL_36_DFFSR_241 gnd vdd FILL
XFILL_36_DFFSR_252 gnd vdd FILL
XFILL_27_3_1 gnd vdd FILL
XFILL_2_3_1 gnd vdd FILL
XFILL_36_DFFSR_263 gnd vdd FILL
XFILL_2_MUX2X1_10 gnd vdd FILL
XFILL_36_DFFSR_274 gnd vdd FILL
XFILL_2_MUX2X1_21 gnd vdd FILL
XFILL_2_MUX2X1_32 gnd vdd FILL
XFILL_2_MUX2X1_43 gnd vdd FILL
XFILL_63_DFFSR_130 gnd vdd FILL
XFILL_5_AOI21X1_15 gnd vdd FILL
XFILL_2_MUX2X1_54 gnd vdd FILL
XFILL_5_AOI21X1_26 gnd vdd FILL
XFILL_2_MUX2X1_65 gnd vdd FILL
XFILL_63_DFFSR_141 gnd vdd FILL
XFILL_2_MUX2X1_76 gnd vdd FILL
XFILL_5_AOI21X1_37 gnd vdd FILL
XFILL_63_DFFSR_152 gnd vdd FILL
XFILL_2_MUX2X1_87 gnd vdd FILL
XFILL_5_AOI21X1_48 gnd vdd FILL
XFILL_5_AOI21X1_59 gnd vdd FILL
XFILL_63_DFFSR_163 gnd vdd FILL
XFILL_63_DFFSR_174 gnd vdd FILL
XFILL_15_OAI22X1_17 gnd vdd FILL
XFILL_2_MUX2X1_98 gnd vdd FILL
XFILL_15_OAI22X1_28 gnd vdd FILL
XFILL_6_MUX2X1_20 gnd vdd FILL
XFILL_63_DFFSR_185 gnd vdd FILL
XFILL_6_MUX2X1_31 gnd vdd FILL
XFILL_15_OAI22X1_39 gnd vdd FILL
XFILL_63_DFFSR_196 gnd vdd FILL
XFILL_6_MUX2X1_42 gnd vdd FILL
XFILL_6_MUX2X1_53 gnd vdd FILL
XFILL_8_NOR2X1_103 gnd vdd FILL
XFILL_11_NAND3X1_9 gnd vdd FILL
XFILL_14_DFFSR_209 gnd vdd FILL
XFILL_8_NOR2X1_114 gnd vdd FILL
XFILL_8_NOR2X1_125 gnd vdd FILL
XFILL_67_DFFSR_140 gnd vdd FILL
XFILL_6_MUX2X1_64 gnd vdd FILL
XFILL_11_7_2 gnd vdd FILL
XFILL_6_MUX2X1_75 gnd vdd FILL
XFILL_67_DFFSR_151 gnd vdd FILL
XFILL_8_NOR2X1_136 gnd vdd FILL
XFILL_0_BUFX4_4 gnd vdd FILL
XFILL_8_NOR2X1_147 gnd vdd FILL
XFILL_6_MUX2X1_86 gnd vdd FILL
XFILL_10_2_1 gnd vdd FILL
XFILL_67_DFFSR_162 gnd vdd FILL
XFILL_6_MUX2X1_97 gnd vdd FILL
XFILL_8_NOR2X1_158 gnd vdd FILL
XFILL_13_BUFX4_2 gnd vdd FILL
XFILL_67_DFFSR_173 gnd vdd FILL
XFILL_67_DFFSR_184 gnd vdd FILL
XFILL_8_NOR2X1_169 gnd vdd FILL
XFILL_14_NAND3X1_60 gnd vdd FILL
XFILL_67_DFFSR_195 gnd vdd FILL
XFILL_41_DFFSR_109 gnd vdd FILL
XFILL_14_NAND3X1_71 gnd vdd FILL
XFILL_18_DFFSR_208 gnd vdd FILL
XFILL_15_NAND3X1_8 gnd vdd FILL
XFILL_18_DFFSR_219 gnd vdd FILL
XFILL_14_NAND3X1_82 gnd vdd FILL
XFILL_14_NAND3X1_93 gnd vdd FILL
XFILL_1_NAND3X1_101 gnd vdd FILL
XFILL_1_NAND3X1_112 gnd vdd FILL
XFILL_1_NAND3X1_123 gnd vdd FILL
XFILL_45_DFFSR_108 gnd vdd FILL
XFILL_45_DFFSR_119 gnd vdd FILL
XFILL_8_MUX2X1_109 gnd vdd FILL
XFILL_49_DFFSR_107 gnd vdd FILL
XFILL_49_DFFSR_118 gnd vdd FILL
XFILL_22_MUX2X1_40 gnd vdd FILL
XFILL_49_DFFSR_129 gnd vdd FILL
XFILL_22_MUX2X1_51 gnd vdd FILL
XFILL_5_OAI22X1_12 gnd vdd FILL
XFILL_22_MUX2X1_62 gnd vdd FILL
XFILL_22_MUX2X1_73 gnd vdd FILL
XFILL_5_OAI22X1_23 gnd vdd FILL
XFILL_22_MUX2X1_84 gnd vdd FILL
XFILL_5_OAI22X1_34 gnd vdd FILL
XFILL_22_MUX2X1_95 gnd vdd FILL
XFILL_5_OAI22X1_45 gnd vdd FILL
XFILL_9_OAI21X1_14 gnd vdd FILL
XFILL_9_OAI21X1_25 gnd vdd FILL
XFILL_18_3_1 gnd vdd FILL
XFILL_9_OAI21X1_36 gnd vdd FILL
XFILL_9_OAI21X1_47 gnd vdd FILL
XFILL_32_7 gnd vdd FILL
XFILL_61_6_2 gnd vdd FILL
XFILL_60_1_1 gnd vdd FILL
XFILL_2_NOR2X1_203 gnd vdd FILL
XFILL_30_DFFSR_130 gnd vdd FILL
XFILL_30_DFFSR_141 gnd vdd FILL
XFILL_30_DFFSR_152 gnd vdd FILL
XFILL_3_INVX8_2 gnd vdd FILL
XFILL_8_NAND2X1_90 gnd vdd FILL
XFILL_30_DFFSR_163 gnd vdd FILL
XFILL_18_5 gnd vdd FILL
XFILL_30_DFFSR_174 gnd vdd FILL
XFILL_30_DFFSR_185 gnd vdd FILL
XFILL_16_CLKBUF1_10 gnd vdd FILL
XFILL_30_DFFSR_196 gnd vdd FILL
XFILL_16_CLKBUF1_21 gnd vdd FILL
XFILL_16_CLKBUF1_32 gnd vdd FILL
XFILL_34_DFFSR_140 gnd vdd FILL
XFILL_34_DFFSR_151 gnd vdd FILL
XFILL_34_DFFSR_162 gnd vdd FILL
XFILL_11_AOI21X1_40 gnd vdd FILL
XFILL_34_DFFSR_173 gnd vdd FILL
XFILL_34_DFFSR_184 gnd vdd FILL
XFILL_11_AOI21X1_51 gnd vdd FILL
XFILL_34_DFFSR_195 gnd vdd FILL
XFILL_20_DFFSR_2 gnd vdd FILL
XFILL_11_AOI21X1_62 gnd vdd FILL
XFILL_11_AOI21X1_73 gnd vdd FILL
XFILL_38_DFFSR_150 gnd vdd FILL
XFILL_38_DFFSR_161 gnd vdd FILL
XFILL_38_DFFSR_172 gnd vdd FILL
XFILL_2_INVX1_16 gnd vdd FILL
XFILL_38_DFFSR_183 gnd vdd FILL
XFILL_2_INVX1_27 gnd vdd FILL
XFILL_2_INVX1_38 gnd vdd FILL
XFILL_38_DFFSR_194 gnd vdd FILL
XFILL_12_DFFSR_108 gnd vdd FILL
XFILL_30_NOR3X1_30 gnd vdd FILL
XFILL_12_DFFSR_119 gnd vdd FILL
XFILL_3_AND2X2_8 gnd vdd FILL
XFILL_2_INVX1_49 gnd vdd FILL
XFILL_30_NOR3X1_41 gnd vdd FILL
XFILL_30_NOR3X1_52 gnd vdd FILL
XFILL_48_DFFSR_19 gnd vdd FILL
XFILL_80_DFFSR_230 gnd vdd FILL
XFILL_80_DFFSR_241 gnd vdd FILL
XFILL_80_DFFSR_252 gnd vdd FILL
XFILL_80_DFFSR_263 gnd vdd FILL
XFILL_80_DFFSR_274 gnd vdd FILL
XFILL_16_DFFSR_107 gnd vdd FILL
XFILL_16_DFFSR_118 gnd vdd FILL
XFILL_16_DFFSR_129 gnd vdd FILL
XFILL_11_AOI21X1_3 gnd vdd FILL
XFILL_0_BUFX4_14 gnd vdd FILL
XFILL_42_DFFSR_6 gnd vdd FILL
XFILL_0_BUFX4_25 gnd vdd FILL
XFILL_84_DFFSR_240 gnd vdd FILL
XFILL_84_DFFSR_251 gnd vdd FILL
XFILL_0_BUFX4_36 gnd vdd FILL
XFILL_84_DFFSR_262 gnd vdd FILL
XFILL_0_BUFX4_47 gnd vdd FILL
XFILL_17_DFFSR_18 gnd vdd FILL
XFILL_17_DFFSR_29 gnd vdd FILL
XFILL_84_DFFSR_273 gnd vdd FILL
XFILL_0_BUFX4_58 gnd vdd FILL
XFILL_0_BUFX4_69 gnd vdd FILL
XFILL_14_MUX2X1_101 gnd vdd FILL
XFILL_14_MUX2X1_112 gnd vdd FILL
XFILL_14_MUX2X1_123 gnd vdd FILL
XFILL_52_6_2 gnd vdd FILL
XFILL_15_AOI21X1_2 gnd vdd FILL
XFILL_14_MUX2X1_134 gnd vdd FILL
XFILL_14_MUX2X1_145 gnd vdd FILL
XFILL_51_1_1 gnd vdd FILL
XFILL_0_INVX1_190 gnd vdd FILL
XFILL_14_MUX2X1_156 gnd vdd FILL
XFILL_57_DFFSR_17 gnd vdd FILL
XFILL_14_MUX2X1_167 gnd vdd FILL
XFILL_12_NOR3X1_19 gnd vdd FILL
XFILL_57_DFFSR_28 gnd vdd FILL
XFILL_14_MUX2X1_178 gnd vdd FILL
XFILL_14_MUX2X1_189 gnd vdd FILL
XFILL_57_DFFSR_39 gnd vdd FILL
XFILL_62_DFFSR_208 gnd vdd FILL
XFILL_62_DFFSR_219 gnd vdd FILL
XFILL_15_OAI21X1_50 gnd vdd FILL
XFILL_16_NOR3X1_18 gnd vdd FILL
XFILL_16_NOR3X1_29 gnd vdd FILL
XFILL_66_DFFSR_207 gnd vdd FILL
XFILL_26_DFFSR_16 gnd vdd FILL
XFILL_66_DFFSR_218 gnd vdd FILL
XFILL_26_DFFSR_27 gnd vdd FILL
XFILL_66_DFFSR_229 gnd vdd FILL
XFILL_26_DFFSR_38 gnd vdd FILL
XFILL_26_DFFSR_49 gnd vdd FILL
XFILL_66_DFFSR_15 gnd vdd FILL
XFILL_66_DFFSR_26 gnd vdd FILL
XFILL_66_DFFSR_37 gnd vdd FILL
XFILL_66_DFFSR_48 gnd vdd FILL
XFILL_66_DFFSR_59 gnd vdd FILL
XNAND3X1_14 INVX1_20/A BUFX4_5/Y NOR2X1_31/Y gnd NAND3X1_16/B vdd NAND3X1
XFILL_21_MUX2X1_180 gnd vdd FILL
XNAND3X1_25 DFFSR_106/Q BUFX4_2/Y NOR2X1_29/Y gnd OAI21X1_32/C vdd NAND3X1
XFILL_21_MUX2X1_191 gnd vdd FILL
XFILL_59_2_1 gnd vdd FILL
XFILL_4_MUX2X1_140 gnd vdd FILL
XNAND3X1_36 INVX2_5/A OAI21X1_43/Y NAND3X1_36/C gnd NAND3X1_43/B vdd NAND3X1
XNAND3X1_47 NOR2X1_33/Y NOR2X1_39/Y NOR3X1_23/Y gnd NOR3X1_3/C vdd NAND3X1
XFILL_4_MUX2X1_151 gnd vdd FILL
XFILL_4_MUX2X1_162 gnd vdd FILL
XNAND3X1_58 BUFX4_57/Y AND2X2_3/B NOR2X1_42/Y gnd OAI22X1_8/D vdd NAND3X1
XFILL_9_DFFSR_17 gnd vdd FILL
XFILL_4_BUFX4_5 gnd vdd FILL
XNAND3X1_69 INVX1_159/A BUFX4_90/Y NOR3X1_51/Y gnd OAI21X1_2/C vdd NAND3X1
XFILL_9_DFFSR_28 gnd vdd FILL
XFILL_7_NAND3X1_106 gnd vdd FILL
XFILL_4_MUX2X1_173 gnd vdd FILL
XFILL_35_DFFSR_14 gnd vdd FILL
XFILL_9_DFFSR_39 gnd vdd FILL
XFILL_7_NAND3X1_117 gnd vdd FILL
XFILL_4_MUX2X1_184 gnd vdd FILL
XFILL_7_NAND3X1_128 gnd vdd FILL
XFILL_35_DFFSR_25 gnd vdd FILL
XNOR2X1_14 NOR2X1_7/B INVX1_3/Y gnd NOR2X1_16/B vdd NOR2X1
XFILL_35_DFFSR_36 gnd vdd FILL
XNOR2X1_25 NOR2X1_25/A OR2X2_1/A gnd NOR2X1_26/B vdd NOR2X1
XFILL_35_DFFSR_47 gnd vdd FILL
XFILL_35_DFFSR_58 gnd vdd FILL
XNOR2X1_36 NOR3X1_52/C NOR2X1_44/B gnd NOR2X1_36/Y vdd NOR2X1
XNOR2X1_47 NOR2X1_47/A NOR2X1_98/B gnd NOR2X1_47/Y vdd NOR2X1
XFILL_35_DFFSR_69 gnd vdd FILL
XNOR2X1_58 OAI21X1_5/Y OAI22X1_5/Y gnd NOR2X1_58/Y vdd NOR2X1
XNOR2X1_69 NOR3X1_39/C INVX2_2/Y gnd NOR2X1_69/Y vdd NOR2X1
XFILL_51_DFFSR_240 gnd vdd FILL
XFILL_75_DFFSR_13 gnd vdd FILL
XFILL_51_DFFSR_251 gnd vdd FILL
XFILL_75_DFFSR_24 gnd vdd FILL
XFILL_51_DFFSR_262 gnd vdd FILL
XFILL_43_6_2 gnd vdd FILL
XFILL_75_DFFSR_35 gnd vdd FILL
XFILL_51_DFFSR_273 gnd vdd FILL
XFILL_75_DFFSR_46 gnd vdd FILL
XFILL_18_MUX2X1_3 gnd vdd FILL
XFILL_75_DFFSR_57 gnd vdd FILL
XFILL_42_1_1 gnd vdd FILL
XFILL_75_DFFSR_68 gnd vdd FILL
XFILL_75_DFFSR_79 gnd vdd FILL
XFILL_3_INVX1_9 gnd vdd FILL
XFILL_55_DFFSR_250 gnd vdd FILL
XFILL_55_DFFSR_261 gnd vdd FILL
XFILL_11_NAND3X1_130 gnd vdd FILL
XFILL_10_CLKBUF1_2 gnd vdd FILL
XFILL_55_DFFSR_272 gnd vdd FILL
XFILL_10_NAND2X1_17 gnd vdd FILL
XFILL_10_NAND2X1_28 gnd vdd FILL
XFILL_44_DFFSR_12 gnd vdd FILL
XFILL_10_NAND2X1_39 gnd vdd FILL
XFILL_0_BUFX2_1 gnd vdd FILL
XFILL_44_DFFSR_23 gnd vdd FILL
XFILL_9_BUFX4_80 gnd vdd FILL
XFILL_44_DFFSR_34 gnd vdd FILL
XFILL_9_BUFX4_91 gnd vdd FILL
XFILL_15_NOR3X1_9 gnd vdd FILL
XFILL_44_DFFSR_45 gnd vdd FILL
XFILL_44_DFFSR_56 gnd vdd FILL
XFILL_82_DFFSR_150 gnd vdd FILL
XFILL_82_DFFSR_161 gnd vdd FILL
XFILL_44_DFFSR_67 gnd vdd FILL
XFILL_59_DFFSR_260 gnd vdd FILL
XFILL_59_DFFSR_271 gnd vdd FILL
XFILL_44_DFFSR_78 gnd vdd FILL
XFILL_14_CLKBUF1_1 gnd vdd FILL
XFILL_82_DFFSR_172 gnd vdd FILL
XFILL_44_DFFSR_89 gnd vdd FILL
XFILL_82_DFFSR_183 gnd vdd FILL
XFILL_82_DFFSR_194 gnd vdd FILL
XFILL_33_DFFSR_207 gnd vdd FILL
XFILL_84_DFFSR_11 gnd vdd FILL
XFILL_2_DFFSR_220 gnd vdd FILL
XFILL_84_DFFSR_22 gnd vdd FILL
XFILL_7_NAND3X1_10 gnd vdd FILL
XFILL_7_NAND3X1_21 gnd vdd FILL
XFILL_33_DFFSR_218 gnd vdd FILL
XFILL_84_DFFSR_33 gnd vdd FILL
XFILL_2_DFFSR_231 gnd vdd FILL
XFILL_2_DFFSR_242 gnd vdd FILL
XFILL_7_NAND3X1_32 gnd vdd FILL
XFILL_33_DFFSR_229 gnd vdd FILL
XFILL_84_DFFSR_44 gnd vdd FILL
XFILL_2_NAND3X1_102 gnd vdd FILL
XFILL_2_DFFSR_253 gnd vdd FILL
XFILL_84_DFFSR_55 gnd vdd FILL
XFILL_2_NAND3X1_113 gnd vdd FILL
XFILL_13_DFFSR_11 gnd vdd FILL
XFILL_2_DFFSR_264 gnd vdd FILL
XFILL_7_NAND3X1_43 gnd vdd FILL
XFILL_86_DFFSR_160 gnd vdd FILL
XFILL_13_DFFSR_22 gnd vdd FILL
XFILL_84_DFFSR_66 gnd vdd FILL
XFILL_2_NAND3X1_124 gnd vdd FILL
XFILL_7_NAND3X1_54 gnd vdd FILL
XFILL_2_DFFSR_275 gnd vdd FILL
XFILL_84_DFFSR_77 gnd vdd FILL
XFILL_7_NAND3X1_65 gnd vdd FILL
XFILL_13_DFFSR_33 gnd vdd FILL
XFILL_86_DFFSR_171 gnd vdd FILL
XFILL_7_NAND3X1_76 gnd vdd FILL
XFILL_84_DFFSR_88 gnd vdd FILL
XFILL_86_DFFSR_182 gnd vdd FILL
XFILL_13_DFFSR_44 gnd vdd FILL
XFILL_84_DFFSR_99 gnd vdd FILL
XFILL_7_NAND3X1_87 gnd vdd FILL
XFILL_86_DFFSR_193 gnd vdd FILL
XFILL_37_DFFSR_206 gnd vdd FILL
XFILL_60_DFFSR_107 gnd vdd FILL
XFILL_13_DFFSR_55 gnd vdd FILL
XFILL_37_DFFSR_217 gnd vdd FILL
XFILL_13_DFFSR_66 gnd vdd FILL
XFILL_60_DFFSR_118 gnd vdd FILL
XFILL_7_NAND3X1_98 gnd vdd FILL
XFILL_13_DFFSR_77 gnd vdd FILL
XFILL_6_DFFSR_230 gnd vdd FILL
XFILL_60_DFFSR_129 gnd vdd FILL
XFILL_6_DFFSR_241 gnd vdd FILL
XFILL_37_DFFSR_228 gnd vdd FILL
XFILL_13_DFFSR_88 gnd vdd FILL
XFILL_13_DFFSR_99 gnd vdd FILL
XFILL_37_DFFSR_239 gnd vdd FILL
XFILL_6_DFFSR_252 gnd vdd FILL
XFILL_7_INVX8_3 gnd vdd FILL
XFILL_53_DFFSR_10 gnd vdd FILL
XFILL_6_DFFSR_263 gnd vdd FILL
XFILL_53_DFFSR_21 gnd vdd FILL
XFILL_6_DFFSR_274 gnd vdd FILL
XFILL_53_DFFSR_32 gnd vdd FILL
XFILL_53_DFFSR_43 gnd vdd FILL
XFILL_3_MUX2X1_19 gnd vdd FILL
XFILL_24_NOR3X1_7 gnd vdd FILL
XFILL_53_DFFSR_54 gnd vdd FILL
XFILL_64_DFFSR_106 gnd vdd FILL
XFILL_53_DFFSR_65 gnd vdd FILL
XFILL_64_DFFSR_117 gnd vdd FILL
XFILL_53_DFFSR_76 gnd vdd FILL
XFILL_64_DFFSR_128 gnd vdd FILL
XFILL_53_DFFSR_87 gnd vdd FILL
XFILL_64_DFFSR_139 gnd vdd FILL
XFILL_53_DFFSR_98 gnd vdd FILL
XFILL_14_AOI21X1_17 gnd vdd FILL
XMUX2X1_10 BUFX4_77/Y INVX1_23/Y MUX2X1_9/S gnd DFFSR_39/D vdd MUX2X1
XFILL_0_NAND2X1_12 gnd vdd FILL
XFILL_14_AOI21X1_28 gnd vdd FILL
XMUX2X1_21 BUFX4_63/Y INVX1_34/Y MUX2X1_22/S gnd DFFSR_3/D vdd MUX2X1
XFILL_0_NAND2X1_23 gnd vdd FILL
XFILL_14_AOI21X1_39 gnd vdd FILL
XFILL_7_MUX2X1_18 gnd vdd FILL
XMUX2X1_32 BUFX4_86/Y INVX1_45/Y NOR2X1_20/Y gnd MUX2X1_32/Y vdd MUX2X1
XFILL_0_NAND2X1_34 gnd vdd FILL
XFILL_24_DFFSR_3 gnd vdd FILL
XNOR2X1_104 OAI21X1_28/Y OAI21X1_27/Y gnd NOR2X1_104/Y vdd NOR2X1
XFILL_7_MUX2X1_29 gnd vdd FILL
XFILL_0_NAND2X1_45 gnd vdd FILL
XMUX2X1_43 INVX1_56/Y BUFX4_77/Y NAND2X1_6/Y gnd MUX2X1_43/Y vdd MUX2X1
XFILL_68_DFFSR_105 gnd vdd FILL
XMUX2X1_54 NOR3X1_1/A BUFX4_83/Y NAND2X1_9/Y gnd MUX2X1_54/Y vdd MUX2X1
XNOR2X1_115 NOR2X1_24/A OAI21X1_46/B gnd AND2X2_8/B vdd NOR2X1
XFILL_0_NAND2X1_56 gnd vdd FILL
XFILL_81_DFFSR_4 gnd vdd FILL
XNOR2X1_126 DFFSR_150/Q AOI21X1_3/B gnd AOI21X1_2/C vdd NOR2X1
XFILL_22_DFFSR_20 gnd vdd FILL
XFILL_68_DFFSR_116 gnd vdd FILL
XMUX2X1_65 MUX2X1_6/B INVX1_78/Y NOR2X1_23/Y gnd MUX2X1_65/Y vdd MUX2X1
XFILL_0_NAND2X1_67 gnd vdd FILL
XFILL_68_DFFSR_127 gnd vdd FILL
XFILL_22_DFFSR_31 gnd vdd FILL
XNOR2X1_137 NOR2X1_138/A INVX1_163/Y gnd INVX1_3/A vdd NOR2X1
XFILL_68_DFFSR_138 gnd vdd FILL
XMUX2X1_76 BUFX4_86/Y INVX1_89/Y NOR2X1_26/B gnd MUX2X1_76/Y vdd MUX2X1
XFILL_0_NAND2X1_78 gnd vdd FILL
XFILL_22_DFFSR_42 gnd vdd FILL
XMUX2X1_87 MUX2X1_87/A BUFX4_86/Y MUX2X1_91/S gnd MUX2X1_87/Y vdd MUX2X1
XFILL_68_DFFSR_149 gnd vdd FILL
XFILL_34_6_2 gnd vdd FILL
XFILL_22_DFFSR_53 gnd vdd FILL
XFILL_0_NAND2X1_89 gnd vdd FILL
XNOR2X1_148 NAND2X1_3/Y INVX1_68/Y gnd NOR2X1_153/B vdd NOR2X1
XNOR2X1_159 DFFSR_82/Q NOR2X1_161/B gnd NOR2X1_159/Y vdd NOR2X1
XFILL_11_OAI21X1_6 gnd vdd FILL
XFILL_22_DFFSR_64 gnd vdd FILL
XMUX2X1_98 MUX2X1_98/A BUFX4_75/Y MUX2X1_99/S gnd DFFSR_79/D vdd MUX2X1
XFILL_0_INVX2_1 gnd vdd FILL
XFILL_33_1_1 gnd vdd FILL
XFILL_22_DFFSR_75 gnd vdd FILL
XFILL_22_DFFSR_86 gnd vdd FILL
XFILL_23_3 gnd vdd FILL
XFILL_22_DFFSR_97 gnd vdd FILL
XFILL_7_NOR3X1_8 gnd vdd FILL
XFILL_62_DFFSR_30 gnd vdd FILL
XFILL_3_AOI22X1_2 gnd vdd FILL
XFILL_62_DFFSR_41 gnd vdd FILL
XFILL_16_2 gnd vdd FILL
XFILL_15_OAI21X1_5 gnd vdd FILL
XFILL_62_DFFSR_52 gnd vdd FILL
XFILL_62_DFFSR_63 gnd vdd FILL
XFILL_62_DFFSR_74 gnd vdd FILL
XFILL_22_DFFSR_250 gnd vdd FILL
XFILL_22_DFFSR_261 gnd vdd FILL
XFILL_62_DFFSR_85 gnd vdd FILL
XFILL_22_DFFSR_272 gnd vdd FILL
XFILL_62_DFFSR_96 gnd vdd FILL
XFILL_3_INVX1_201 gnd vdd FILL
XFILL_3_INVX1_212 gnd vdd FILL
XFILL_26_CLKBUF1_11 gnd vdd FILL
XFILL_5_DFFSR_10 gnd vdd FILL
XFILL_26_CLKBUF1_22 gnd vdd FILL
XFILL_3_INVX1_223 gnd vdd FILL
XDFFSR_2 DFFSR_2/Q DFFSR_2/CLK DFFSR_2/R vdd DFFSR_2/D gnd vdd DFFSR
XFILL_5_DFFSR_21 gnd vdd FILL
XFILL_26_CLKBUF1_33 gnd vdd FILL
XFILL_7_AOI22X1_1 gnd vdd FILL
XFILL_5_DFFSR_32 gnd vdd FILL
XFILL_5_DFFSR_43 gnd vdd FILL
XFILL_5_DFFSR_54 gnd vdd FILL
XFILL_46_DFFSR_7 gnd vdd FILL
XFILL_0_AOI22X1_10 gnd vdd FILL
XFILL_5_DFFSR_65 gnd vdd FILL
XFILL_26_DFFSR_260 gnd vdd FILL
XFILL_26_DFFSR_271 gnd vdd FILL
XFILL_31_DFFSR_40 gnd vdd FILL
XFILL_9_CLKBUF1_15 gnd vdd FILL
XFILL_5_DFFSR_76 gnd vdd FILL
XFILL_31_DFFSR_51 gnd vdd FILL
XFILL_7_INVX1_200 gnd vdd FILL
XFILL_23_MUX2X1_16 gnd vdd FILL
XFILL_5_DFFSR_87 gnd vdd FILL
XFILL_31_DFFSR_62 gnd vdd FILL
XFILL_9_CLKBUF1_26 gnd vdd FILL
XFILL_7_INVX1_211 gnd vdd FILL
XFILL_5_DFFSR_98 gnd vdd FILL
XFILL_31_DFFSR_73 gnd vdd FILL
XFILL_23_MUX2X1_27 gnd vdd FILL
XFILL_9_CLKBUF1_37 gnd vdd FILL
XFILL_7_INVX1_222 gnd vdd FILL
XFILL_31_DFFSR_84 gnd vdd FILL
XFILL_4_AOI21X1_12 gnd vdd FILL
XFILL_23_MUX2X1_38 gnd vdd FILL
XFILL_14_10 gnd vdd FILL
XFILL_23_MUX2X1_49 gnd vdd FILL
XFILL_31_DFFSR_95 gnd vdd FILL
XFILL_4_AOI21X1_23 gnd vdd FILL
XFILL_4_AOI21X1_34 gnd vdd FILL
XFILL_4_AOI21X1_45 gnd vdd FILL
XFILL_53_DFFSR_160 gnd vdd FILL
XFILL_4_AOI21X1_56 gnd vdd FILL
XFILL_4_AOI21X1_67 gnd vdd FILL
XFILL_14_OAI22X1_14 gnd vdd FILL
XFILL_53_DFFSR_171 gnd vdd FILL
XFILL_14_OAI22X1_25 gnd vdd FILL
XFILL_53_DFFSR_182 gnd vdd FILL
XFILL_71_DFFSR_50 gnd vdd FILL
XFILL_4_AOI21X1_78 gnd vdd FILL
XFILL_53_DFFSR_193 gnd vdd FILL
XFILL_14_OAI22X1_36 gnd vdd FILL
XFILL_71_DFFSR_61 gnd vdd FILL
XFILL_14_OAI22X1_47 gnd vdd FILL
XINVX1_17 INVX1_17/A gnd MUX2X1_4/A vdd INVX1
XFILL_7_NOR2X1_100 gnd vdd FILL
XFILL_71_DFFSR_72 gnd vdd FILL
XFILL_71_DFFSR_83 gnd vdd FILL
XINVX1_28 INVX1_28/A gnd INVX1_28/Y vdd INVX1
XFILL_7_NOR2X1_111 gnd vdd FILL
XFILL_71_DFFSR_94 gnd vdd FILL
XFILL_7_NOR2X1_122 gnd vdd FILL
XINVX1_39 INVX1_39/A gnd INVX1_39/Y vdd INVX1
XFILL_7_NOR2X1_133 gnd vdd FILL
XFILL_7_NOR2X1_144 gnd vdd FILL
XFILL_7_NOR2X1_155 gnd vdd FILL
XFILL_57_DFFSR_170 gnd vdd FILL
XFILL_7_NOR2X1_166 gnd vdd FILL
XFILL_57_DFFSR_181 gnd vdd FILL
XFILL_7_NOR2X1_177 gnd vdd FILL
XFILL_57_DFFSR_192 gnd vdd FILL
XFILL_31_DFFSR_106 gnd vdd FILL
XFILL_7_NOR2X1_188 gnd vdd FILL
XFILL_0_DFFSR_130 gnd vdd FILL
XFILL_7_NOR2X1_199 gnd vdd FILL
XFILL_11_NOR3X1_2 gnd vdd FILL
XFILL_31_DFFSR_117 gnd vdd FILL
XNAND2X1_80 NOR2X1_105/Y NOR2X1_104/Y gnd NOR3X1_47/C vdd NAND2X1
XFILL_31_DFFSR_128 gnd vdd FILL
XFILL_0_DFFSR_141 gnd vdd FILL
XNAND2X1_91 INVX1_131/A INVX1_133/Y gnd NOR2X1_21/A vdd NAND2X1
XFILL_31_DFFSR_139 gnd vdd FILL
XFILL_13_NAND3X1_90 gnd vdd FILL
XFILL_0_DFFSR_152 gnd vdd FILL
XFILL_40_DFFSR_60 gnd vdd FILL
XFILL_11_NOR2X1_205 gnd vdd FILL
XFILL_0_DFFSR_163 gnd vdd FILL
XFILL_40_DFFSR_71 gnd vdd FILL
XFILL_40_DFFSR_82 gnd vdd FILL
XFILL_0_DFFSR_174 gnd vdd FILL
XFILL_40_DFFSR_93 gnd vdd FILL
XFILL_0_DFFSR_185 gnd vdd FILL
XFILL_0_DFFSR_196 gnd vdd FILL
XFILL_25_6_2 gnd vdd FILL
XFILL_35_DFFSR_105 gnd vdd FILL
XFILL_0_6_2 gnd vdd FILL
XFILL_35_DFFSR_116 gnd vdd FILL
XFILL_4_DFFSR_140 gnd vdd FILL
XFILL_35_DFFSR_127 gnd vdd FILL
XFILL_24_1_1 gnd vdd FILL
XFILL_35_DFFSR_138 gnd vdd FILL
XFILL_4_DFFSR_151 gnd vdd FILL
XFILL_35_DFFSR_149 gnd vdd FILL
XFILL_4_DFFSR_162 gnd vdd FILL
XFILL_80_DFFSR_70 gnd vdd FILL
XFILL_4_DFFSR_173 gnd vdd FILL
XFILL_80_DFFSR_81 gnd vdd FILL
XFILL_4_DFFSR_184 gnd vdd FILL
XFILL_80_DFFSR_92 gnd vdd FILL
XFILL_4_DFFSR_195 gnd vdd FILL
XFILL_39_DFFSR_104 gnd vdd FILL
XFILL_7_MUX2X1_106 gnd vdd FILL
XFILL_7_MUX2X1_117 gnd vdd FILL
XFILL_39_DFFSR_115 gnd vdd FILL
XFILL_39_DFFSR_126 gnd vdd FILL
XFILL_7_MUX2X1_128 gnd vdd FILL
XFILL_39_DFFSR_137 gnd vdd FILL
XFILL_8_DFFSR_150 gnd vdd FILL
XFILL_7_MUX2X1_139 gnd vdd FILL
XFILL_8_DFFSR_161 gnd vdd FILL
XFILL_39_DFFSR_148 gnd vdd FILL
XFILL_8_BUFX4_6 gnd vdd FILL
XFILL_4_OAI22X1_20 gnd vdd FILL
XFILL_8_DFFSR_172 gnd vdd FILL
XFILL_12_MUX2X1_70 gnd vdd FILL
XFILL_39_DFFSR_159 gnd vdd FILL
XFILL_12_MUX2X1_81 gnd vdd FILL
XFILL_4_OAI22X1_31 gnd vdd FILL
XFILL_8_DFFSR_183 gnd vdd FILL
XFILL_4_OAI22X1_42 gnd vdd FILL
XFILL_12_MUX2X1_92 gnd vdd FILL
XFILL_31_NOR3X1_17 gnd vdd FILL
XFILL_8_DFFSR_194 gnd vdd FILL
XFILL_0_NOR3X1_30 gnd vdd FILL
XFILL_8_OAI21X1_11 gnd vdd FILL
XFILL_31_NOR3X1_28 gnd vdd FILL
XFILL_0_NOR3X1_41 gnd vdd FILL
XFILL_0_NOR3X1_52 gnd vdd FILL
XFILL_31_NOR3X1_39 gnd vdd FILL
XFILL_8_OAI21X1_22 gnd vdd FILL
XFILL_81_DFFSR_206 gnd vdd FILL
XFILL_8_OAI21X1_33 gnd vdd FILL
XFILL_8_OAI21X1_44 gnd vdd FILL
XFILL_81_DFFSR_217 gnd vdd FILL
XFILL_81_DFFSR_228 gnd vdd FILL
XFILL_81_DFFSR_239 gnd vdd FILL
XFILL_16_MUX2X1_80 gnd vdd FILL
XFILL_16_MUX2X1_91 gnd vdd FILL
XFILL_4_NOR3X1_40 gnd vdd FILL
XFILL_4_NOR3X1_51 gnd vdd FILL
XFILL_85_DFFSR_205 gnd vdd FILL
XFILL_1_NOR2X1_200 gnd vdd FILL
XFILL_85_DFFSR_216 gnd vdd FILL
XFILL_85_DFFSR_227 gnd vdd FILL
XFILL_85_DFFSR_238 gnd vdd FILL
XFILL_8_7_2 gnd vdd FILL
XFILL_20_DFFSR_160 gnd vdd FILL
XFILL_85_DFFSR_249 gnd vdd FILL
XFILL_7_2_1 gnd vdd FILL
XFILL_3_NOR3X1_1 gnd vdd FILL
XFILL_20_DFFSR_171 gnd vdd FILL
XFILL_1_INVX1_100 gnd vdd FILL
XFILL_20_DFFSR_182 gnd vdd FILL
XFILL_20_DFFSR_193 gnd vdd FILL
XFILL_1_INVX1_111 gnd vdd FILL
XFILL_8_NOR3X1_50 gnd vdd FILL
XFILL_1_INVX1_122 gnd vdd FILL
XFILL_4_BUFX2_2 gnd vdd FILL
XFILL_1_INVX1_133 gnd vdd FILL
XFILL_1_INVX1_144 gnd vdd FILL
XFILL_15_CLKBUF1_40 gnd vdd FILL
XFILL_1_INVX1_155 gnd vdd FILL
XFILL_1_INVX1_166 gnd vdd FILL
XFILL_8_NAND3X1_107 gnd vdd FILL
XFILL_1_INVX1_177 gnd vdd FILL
XFILL_1_INVX1_188 gnd vdd FILL
XFILL_24_DFFSR_170 gnd vdd FILL
XFILL_8_NAND3X1_118 gnd vdd FILL
XFILL_24_DFFSR_181 gnd vdd FILL
XFILL_1_INVX1_199 gnd vdd FILL
XFILL_5_INVX1_110 gnd vdd FILL
XFILL_8_NAND3X1_129 gnd vdd FILL
XFILL_24_DFFSR_192 gnd vdd FILL
XFILL_5_INVX1_121 gnd vdd FILL
XFILL_10_AOI21X1_70 gnd vdd FILL
XFILL_5_INVX1_132 gnd vdd FILL
XFILL_10_AOI21X1_81 gnd vdd FILL
XFILL_5_INVX1_143 gnd vdd FILL
XFILL_5_INVX1_154 gnd vdd FILL
XFILL_63_DFFSR_1 gnd vdd FILL
XFILL_16_6_2 gnd vdd FILL
XFILL_5_INVX1_165 gnd vdd FILL
XFILL_1_DFFSR_80 gnd vdd FILL
XFILL_5_INVX1_176 gnd vdd FILL
XFILL_5_INVX1_187 gnd vdd FILL
XFILL_15_1_1 gnd vdd FILL
XFILL_28_DFFSR_180 gnd vdd FILL
XFILL_5_INVX1_198 gnd vdd FILL
XFILL_1_DFFSR_91 gnd vdd FILL
XFILL_28_DFFSR_191 gnd vdd FILL
XFILL_70_DFFSR_260 gnd vdd FILL
XFILL_12_NAND3X1_120 gnd vdd FILL
XFILL_12_NAND3X1_131 gnd vdd FILL
XFILL_70_DFFSR_271 gnd vdd FILL
XFILL_3_OAI22X1_5 gnd vdd FILL
XFILL_28_DFFSR_4 gnd vdd FILL
XFILL_74_DFFSR_270 gnd vdd FILL
XFILL_85_DFFSR_5 gnd vdd FILL
XFILL_13_MUX2X1_120 gnd vdd FILL
XFILL_7_OAI22X1_4 gnd vdd FILL
XFILL_4_INVX2_2 gnd vdd FILL
XFILL_3_NAND3X1_103 gnd vdd FILL
XFILL_13_MUX2X1_131 gnd vdd FILL
XFILL_13_MUX2X1_142 gnd vdd FILL
XFILL_13_MUX2X1_153 gnd vdd FILL
XFILL_3_NAND3X1_114 gnd vdd FILL
XFILL_3_NAND3X1_125 gnd vdd FILL
XFILL_13_MUX2X1_164 gnd vdd FILL
XFILL_13_MUX2X1_175 gnd vdd FILL
XFILL_13_MUX2X1_186 gnd vdd FILL
XFILL_52_DFFSR_205 gnd vdd FILL
XFILL_52_DFFSR_216 gnd vdd FILL
XFILL_52_DFFSR_227 gnd vdd FILL
XFILL_52_DFFSR_238 gnd vdd FILL
XFILL_52_DFFSR_249 gnd vdd FILL
XFILL_66_5_2 gnd vdd FILL
XFILL_56_DFFSR_204 gnd vdd FILL
XFILL_65_0_1 gnd vdd FILL
XFILL_56_DFFSR_215 gnd vdd FILL
XFILL_56_DFFSR_226 gnd vdd FILL
XFILL_56_DFFSR_237 gnd vdd FILL
XFILL_56_DFFSR_248 gnd vdd FILL
XFILL_56_DFFSR_259 gnd vdd FILL
XFILL_83_DFFSR_104 gnd vdd FILL
XFILL_83_DFFSR_115 gnd vdd FILL
XFILL_83_DFFSR_126 gnd vdd FILL
XFILL_83_DFFSR_137 gnd vdd FILL
XFILL_83_DFFSR_148 gnd vdd FILL
XFILL_83_DFFSR_159 gnd vdd FILL
XFILL_3_DFFSR_207 gnd vdd FILL
XFILL_87_DFFSR_103 gnd vdd FILL
XFILL_0_NAND3X1_7 gnd vdd FILL
XFILL_87_DFFSR_114 gnd vdd FILL
XFILL_3_DFFSR_218 gnd vdd FILL
XFILL_3_DFFSR_229 gnd vdd FILL
XFILL_87_DFFSR_125 gnd vdd FILL
XFILL_87_DFFSR_136 gnd vdd FILL
XFILL_14_BUFX4_30 gnd vdd FILL
XFILL_87_DFFSR_147 gnd vdd FILL
XFILL_87_DFFSR_158 gnd vdd FILL
XFILL_14_BUFX4_41 gnd vdd FILL
XFILL_3_MUX2X1_170 gnd vdd FILL
XFILL_11_BUFX4_105 gnd vdd FILL
XFILL_14_BUFX4_52 gnd vdd FILL
XFILL_87_DFFSR_169 gnd vdd FILL
XFILL_3_MUX2X1_181 gnd vdd FILL
XFILL_19_CLKBUF1_9 gnd vdd FILL
XFILL_14_BUFX4_63 gnd vdd FILL
XFILL_3_MUX2X1_192 gnd vdd FILL
XFILL_7_DFFSR_206 gnd vdd FILL
XDFFSR_220 INVX1_78/A DFFSR_47/CLK DFFSR_26/R vdd MUX2X1_65/Y gnd vdd DFFSR
XFILL_14_BUFX4_74 gnd vdd FILL
XFILL_14_BUFX4_85 gnd vdd FILL
XFILL_7_DFFSR_217 gnd vdd FILL
XFILL_4_NAND3X1_6 gnd vdd FILL
XDFFSR_231 INVX1_63/A CLKBUF1_26/Y DFFSR_25/R vdd MUX2X1_50/Y gnd vdd DFFSR
XFILL_14_BUFX4_96 gnd vdd FILL
XDFFSR_242 INVX1_56/A CLKBUF1_34/Y BUFX4_23/Y vdd MUX2X1_43/Y gnd vdd DFFSR
XFILL_7_DFFSR_228 gnd vdd FILL
XDFFSR_253 NOR2X1_18/A DFFSR_6/CLK BUFX4_54/Y vdd DFFSR_253/D gnd vdd DFFSR
XFILL_7_DFFSR_239 gnd vdd FILL
XDFFSR_264 INVX1_40/A DFFSR_1/CLK BUFX4_54/Y vdd MUX2X1_27/Y gnd vdd DFFSR
XDFFSR_275 DFFSR_275/Q DFFSR_9/CLK DFFSR_9/R vdd DFFSR_275/D gnd vdd DFFSR
XFILL_15_BUFX4_104 gnd vdd FILL
XFILL_63_DFFSR_19 gnd vdd FILL
XFILL_41_DFFSR_270 gnd vdd FILL
XFILL_8_NAND3X1_5 gnd vdd FILL
XFILL_32_DFFSR_18 gnd vdd FILL
XFILL_32_DFFSR_29 gnd vdd FILL
XFILL_9_AND2X2_1 gnd vdd FILL
XFILL_57_5_2 gnd vdd FILL
XFILL_7_OAI22X1_19 gnd vdd FILL
XFILL_56_0_1 gnd vdd FILL
XFILL_72_DFFSR_180 gnd vdd FILL
XFILL_72_DFFSR_17 gnd vdd FILL
XFILL_72_DFFSR_191 gnd vdd FILL
XFILL_72_DFFSR_28 gnd vdd FILL
XFILL_23_DFFSR_204 gnd vdd FILL
XFILL_23_DFFSR_215 gnd vdd FILL
XFILL_72_DFFSR_39 gnd vdd FILL
XFILL_23_DFFSR_226 gnd vdd FILL
XFILL_15_MUX2X1_7 gnd vdd FILL
XFILL_23_DFFSR_237 gnd vdd FILL
XFILL_6_NAND3X1_40 gnd vdd FILL
XFILL_23_DFFSR_248 gnd vdd FILL
XFILL_6_NAND3X1_51 gnd vdd FILL
XFILL_23_DFFSR_259 gnd vdd FILL
XFILL_6_NAND3X1_62 gnd vdd FILL
XFILL_6_NAND3X1_73 gnd vdd FILL
XFILL_6_NAND3X1_84 gnd vdd FILL
XFILL_76_DFFSR_190 gnd vdd FILL
XFILL_50_DFFSR_104 gnd vdd FILL
XFILL_6_NAND3X1_95 gnd vdd FILL
XFILL_27_DFFSR_203 gnd vdd FILL
XFILL_6_BUFX4_40 gnd vdd FILL
XFILL_50_DFFSR_115 gnd vdd FILL
XFILL_27_DFFSR_214 gnd vdd FILL
XFILL_6_BUFX4_51 gnd vdd FILL
XFILL_50_DFFSR_126 gnd vdd FILL
XFILL_50_DFFSR_137 gnd vdd FILL
XFILL_27_DFFSR_225 gnd vdd FILL
XFILL_40_4_2 gnd vdd FILL
XFILL_41_DFFSR_16 gnd vdd FILL
XFILL_27_DFFSR_236 gnd vdd FILL
XFILL_6_BUFX4_62 gnd vdd FILL
XFILL_50_DFFSR_148 gnd vdd FILL
XFILL_6_BUFX4_73 gnd vdd FILL
XFILL_27_DFFSR_247 gnd vdd FILL
XFILL_41_DFFSR_27 gnd vdd FILL
XFILL_6_BUFX4_84 gnd vdd FILL
XFILL_41_DFFSR_38 gnd vdd FILL
XFILL_27_DFFSR_258 gnd vdd FILL
XFILL_50_DFFSR_159 gnd vdd FILL
XFILL_6_BUFX4_95 gnd vdd FILL
XFILL_27_DFFSR_269 gnd vdd FILL
XFILL_41_DFFSR_49 gnd vdd FILL
XFILL_54_DFFSR_103 gnd vdd FILL
XFILL_8_BUFX2_3 gnd vdd FILL
XFILL_54_DFFSR_114 gnd vdd FILL
XFILL_18_CLKBUF1_17 gnd vdd FILL
XFILL_18_CLKBUF1_28 gnd vdd FILL
XFILL_54_DFFSR_125 gnd vdd FILL
XFILL_54_DFFSR_136 gnd vdd FILL
XFILL_18_CLKBUF1_39 gnd vdd FILL
XFILL_81_DFFSR_15 gnd vdd FILL
XFILL_54_DFFSR_147 gnd vdd FILL
XFILL_13_AOI21X1_14 gnd vdd FILL
XFILL_81_DFFSR_26 gnd vdd FILL
XFILL_54_DFFSR_158 gnd vdd FILL
XFILL_81_DFFSR_37 gnd vdd FILL
XFILL_13_AOI21X1_25 gnd vdd FILL
XFILL_13_AOI21X1_36 gnd vdd FILL
XFILL_54_DFFSR_169 gnd vdd FILL
XFILL_81_DFFSR_48 gnd vdd FILL
XFILL_13_AOI21X1_47 gnd vdd FILL
XFILL_58_DFFSR_102 gnd vdd FILL
XFILL_10_DFFSR_15 gnd vdd FILL
XFILL_81_DFFSR_59 gnd vdd FILL
XFILL_10_DFFSR_26 gnd vdd FILL
XFILL_13_AOI21X1_58 gnd vdd FILL
XFILL_13_AOI21X1_69 gnd vdd FILL
XFILL_10_DFFSR_37 gnd vdd FILL
XFILL_58_DFFSR_113 gnd vdd FILL
XFILL_58_DFFSR_124 gnd vdd FILL
XFILL_10_DFFSR_48 gnd vdd FILL
XFILL_58_DFFSR_135 gnd vdd FILL
XFILL_67_DFFSR_2 gnd vdd FILL
XFILL_58_DFFSR_146 gnd vdd FILL
XFILL_10_DFFSR_59 gnd vdd FILL
XFILL_58_DFFSR_157 gnd vdd FILL
XFILL_8_NOR2X1_8 gnd vdd FILL
XFILL_58_DFFSR_168 gnd vdd FILL
XFILL_58_DFFSR_179 gnd vdd FILL
XFILL_1_DFFSR_106 gnd vdd FILL
XFILL_50_DFFSR_14 gnd vdd FILL
XFILL_1_DFFSR_117 gnd vdd FILL
XFILL_50_DFFSR_25 gnd vdd FILL
XFILL_50_DFFSR_36 gnd vdd FILL
XFILL_1_DFFSR_128 gnd vdd FILL
XFILL_1_DFFSR_139 gnd vdd FILL
XFILL_50_DFFSR_47 gnd vdd FILL
XFILL_50_DFFSR_58 gnd vdd FILL
XFILL_50_DFFSR_69 gnd vdd FILL
XFILL_5_DFFSR_105 gnd vdd FILL
XFILL_48_5_2 gnd vdd FILL
XFILL_5_DFFSR_116 gnd vdd FILL
XFILL_7_MUX2X1_6 gnd vdd FILL
XFILL_5_DFFSR_127 gnd vdd FILL
XFILL_5_DFFSR_138 gnd vdd FILL
XFILL_25_CLKBUF1_30 gnd vdd FILL
XFILL_5_DFFSR_149 gnd vdd FILL
XFILL_47_0_1 gnd vdd FILL
XFILL_0_AOI21X1_1 gnd vdd FILL
XFILL_25_CLKBUF1_41 gnd vdd FILL
XFILL_51_DFFSR_8 gnd vdd FILL
XFILL_9_NAND3X1_108 gnd vdd FILL
XFILL_8_CLKBUF1_12 gnd vdd FILL
XFILL_9_DFFSR_104 gnd vdd FILL
XFILL_8_CLKBUF1_23 gnd vdd FILL
XFILL_9_NAND3X1_119 gnd vdd FILL
XFILL_13_MUX2X1_13 gnd vdd FILL
XFILL_9_DFFSR_115 gnd vdd FILL
XFILL_8_CLKBUF1_34 gnd vdd FILL
XFILL_9_DFFSR_126 gnd vdd FILL
XFILL_13_MUX2X1_24 gnd vdd FILL
XFILL_9_DFFSR_137 gnd vdd FILL
XFILL_13_MUX2X1_35 gnd vdd FILL
XFILL_3_AOI21X1_20 gnd vdd FILL
XFILL_9_DFFSR_148 gnd vdd FILL
XFILL_16_MUX2X1_108 gnd vdd FILL
XFILL_13_MUX2X1_46 gnd vdd FILL
XFILL_16_MUX2X1_119 gnd vdd FILL
XFILL_9_DFFSR_159 gnd vdd FILL
XFILL_3_AOI21X1_31 gnd vdd FILL
XFILL_13_MUX2X1_57 gnd vdd FILL
XFILL_3_AOI21X1_42 gnd vdd FILL
XFILL_13_MUX2X1_68 gnd vdd FILL
XFILL_13_MUX2X1_79 gnd vdd FILL
XFILL_30_NOR3X1_9 gnd vdd FILL
XFILL_1_NOR3X1_17 gnd vdd FILL
XFILL_3_AOI21X1_53 gnd vdd FILL
XOAI21X1_12 OAI21X1_35/A NOR2X1_20/A BUFX2_9/A gnd OAI21X1_12/Y vdd OAI21X1
XFILL_13_OAI22X1_11 gnd vdd FILL
XFILL_3_AOI21X1_64 gnd vdd FILL
XFILL_1_NOR3X1_28 gnd vdd FILL
XFILL_3_AOI21X1_75 gnd vdd FILL
XOAI21X1_23 NOR3X1_48/B NOR3X1_48/C INVX2_3/Y gnd OAI21X1_23/Y vdd OAI21X1
XFILL_13_OAI22X1_22 gnd vdd FILL
XFILL_17_MUX2X1_12 gnd vdd FILL
XFILL_43_DFFSR_190 gnd vdd FILL
XFILL_1_NOR3X1_39 gnd vdd FILL
XOAI21X1_34 OAI21X1_41/A AOI22X1_3/A INVX2_4/A gnd OAI21X1_34/Y vdd OAI21X1
XFILL_13_OAI22X1_33 gnd vdd FILL
XFILL_31_4_2 gnd vdd FILL
XFILL_17_MUX2X1_23 gnd vdd FILL
XFILL_13_OAI22X1_44 gnd vdd FILL
XOAI21X1_45 OAI21X1_45/A OAI21X1_45/B INVX2_5/A gnd OAI21X1_45/Y vdd OAI21X1
XFILL_17_MUX2X1_34 gnd vdd FILL
XFILL_17_MUX2X1_45 gnd vdd FILL
XFILL_17_MUX2X1_56 gnd vdd FILL
XFILL_2_DFFSR_14 gnd vdd FILL
XFILL_6_NOR2X1_130 gnd vdd FILL
XFILL_6_NOR2X1_141 gnd vdd FILL
XFILL_17_MUX2X1_67 gnd vdd FILL
XFILL_5_NOR3X1_16 gnd vdd FILL
XFILL_17_MUX2X1_78 gnd vdd FILL
XFILL_2_DFFSR_25 gnd vdd FILL
XFILL_6_NOR2X1_152 gnd vdd FILL
XFILL_13_NAND3X1_110 gnd vdd FILL
XFILL_5_NOR3X1_27 gnd vdd FILL
XFILL_2_DFFSR_36 gnd vdd FILL
XFILL_13_NAND3X1_121 gnd vdd FILL
XFILL_17_MUX2X1_89 gnd vdd FILL
XFILL_6_INVX1_1 gnd vdd FILL
XFILL_6_NOR2X1_163 gnd vdd FILL
XFILL_2_DFFSR_47 gnd vdd FILL
XFILL_2_DFFSR_58 gnd vdd FILL
XFILL_5_NOR3X1_38 gnd vdd FILL
XFILL_6_NOR2X1_174 gnd vdd FILL
XFILL_13_NAND3X1_132 gnd vdd FILL
XFILL_5_NOR3X1_49 gnd vdd FILL
XFILL_21_DFFSR_103 gnd vdd FILL
XFILL_2_DFFSR_69 gnd vdd FILL
XFILL_6_NOR2X1_185 gnd vdd FILL
XFILL_21_DFFSR_114 gnd vdd FILL
XFILL_6_NOR2X1_196 gnd vdd FILL
XFILL_21_DFFSR_125 gnd vdd FILL
XFILL_21_DFFSR_136 gnd vdd FILL
XFILL_10_NOR2X1_202 gnd vdd FILL
XFILL_21_DFFSR_147 gnd vdd FILL
XFILL_21_DFFSR_158 gnd vdd FILL
XFILL_9_NOR3X1_15 gnd vdd FILL
XFILL_9_NOR3X1_26 gnd vdd FILL
XFILL_21_DFFSR_169 gnd vdd FILL
XFILL_4_INVX1_90 gnd vdd FILL
XFILL_4_BUFX2_10 gnd vdd FILL
XFILL_9_NOR3X1_37 gnd vdd FILL
XFILL_25_DFFSR_102 gnd vdd FILL
XFILL_2_INVX1_109 gnd vdd FILL
XFILL_9_NOR3X1_48 gnd vdd FILL
XFILL_25_DFFSR_113 gnd vdd FILL
XFILL_25_DFFSR_124 gnd vdd FILL
XFILL_23_MUX2X1_110 gnd vdd FILL
XFILL_25_DFFSR_135 gnd vdd FILL
XFILL_25_DFFSR_146 gnd vdd FILL
XFILL_23_MUX2X1_121 gnd vdd FILL
XFILL_23_MUX2X1_132 gnd vdd FILL
XFILL_4_NAND3X1_104 gnd vdd FILL
XFILL_25_DFFSR_157 gnd vdd FILL
XFILL_23_MUX2X1_143 gnd vdd FILL
XFILL_23_MUX2X1_154 gnd vdd FILL
XFILL_4_NAND3X1_115 gnd vdd FILL
XFILL_25_DFFSR_168 gnd vdd FILL
XFILL_25_DFFSR_179 gnd vdd FILL
XFILL_4_NAND3X1_126 gnd vdd FILL
XFILL_23_MUX2X1_165 gnd vdd FILL
XFILL_6_MUX2X1_103 gnd vdd FILL
XFILL_29_DFFSR_101 gnd vdd FILL
XFILL_6_INVX1_108 gnd vdd FILL
XFILL_6_MUX2X1_114 gnd vdd FILL
XFILL_29_DFFSR_112 gnd vdd FILL
XFILL_23_MUX2X1_176 gnd vdd FILL
XFILL_6_INVX1_119 gnd vdd FILL
XFILL_6_MUX2X1_125 gnd vdd FILL
XFILL_23_MUX2X1_187 gnd vdd FILL
XFILL_29_DFFSR_123 gnd vdd FILL
XFILL_29_DFFSR_134 gnd vdd FILL
XFILL_6_MUX2X1_136 gnd vdd FILL
XFILL_29_DFFSR_145 gnd vdd FILL
XFILL_6_MUX2X1_147 gnd vdd FILL
XFILL_29_DFFSR_156 gnd vdd FILL
XFILL_6_MUX2X1_158 gnd vdd FILL
XFILL_39_5_2 gnd vdd FILL
XFILL_6_MUX2X1_169 gnd vdd FILL
XFILL_29_DFFSR_167 gnd vdd FILL
XFILL_19_DFFSR_70 gnd vdd FILL
XFILL_29_DFFSR_178 gnd vdd FILL
XFILL_21_NOR3X1_14 gnd vdd FILL
XFILL_38_0_1 gnd vdd FILL
XFILL_19_DFFSR_81 gnd vdd FILL
XFILL_19_DFFSR_92 gnd vdd FILL
XFILL_3_OAI22X1_50 gnd vdd FILL
XFILL_29_DFFSR_189 gnd vdd FILL
XFILL_21_NOR3X1_25 gnd vdd FILL
XFILL_21_NOR3X1_36 gnd vdd FILL
XFILL_7_OAI21X1_30 gnd vdd FILL
XFILL_21_NOR3X1_47 gnd vdd FILL
XFILL_71_DFFSR_203 gnd vdd FILL
XFILL_7_OAI21X1_41 gnd vdd FILL
XFILL_71_DFFSR_214 gnd vdd FILL
XFILL_71_DFFSR_225 gnd vdd FILL
XFILL_71_DFFSR_236 gnd vdd FILL
XFILL_71_DFFSR_247 gnd vdd FILL
XFILL_59_DFFSR_80 gnd vdd FILL
XFILL_25_NOR3X1_13 gnd vdd FILL
XFILL_71_DFFSR_258 gnd vdd FILL
XFILL_71_DFFSR_269 gnd vdd FILL
XFILL_25_NOR3X1_24 gnd vdd FILL
XFILL_59_DFFSR_91 gnd vdd FILL
XFILL_25_NOR3X1_35 gnd vdd FILL
XFILL_75_DFFSR_202 gnd vdd FILL
XFILL_25_NOR3X1_46 gnd vdd FILL
XFILL_75_DFFSR_213 gnd vdd FILL
XFILL_4_NOR2X1_1 gnd vdd FILL
XFILL_75_DFFSR_224 gnd vdd FILL
XFILL_50_7_0 gnd vdd FILL
XFILL_75_DFFSR_235 gnd vdd FILL
XFILL_22_4_2 gnd vdd FILL
XFILL_75_DFFSR_246 gnd vdd FILL
XFILL_29_NOR3X1_12 gnd vdd FILL
XFILL_75_DFFSR_257 gnd vdd FILL
XFILL_75_DFFSR_268 gnd vdd FILL
XFILL_29_NOR3X1_23 gnd vdd FILL
XFILL_29_NOR3X1_34 gnd vdd FILL
XFILL_30_CLKBUF1_9 gnd vdd FILL
XFILL_10_DFFSR_190 gnd vdd FILL
XFILL_79_DFFSR_201 gnd vdd FILL
XFILL_29_NOR3X1_45 gnd vdd FILL
XFILL_79_DFFSR_212 gnd vdd FILL
XFILL_28_DFFSR_90 gnd vdd FILL
XFILL_79_DFFSR_223 gnd vdd FILL
XFILL_79_DFFSR_234 gnd vdd FILL
XFILL_79_DFFSR_245 gnd vdd FILL
XFILL_79_DFFSR_256 gnd vdd FILL
XFILL_79_DFFSR_267 gnd vdd FILL
XFILL_34_CLKBUF1_8 gnd vdd FILL
XFILL_11_DFFSR_1 gnd vdd FILL
XFILL_9_NAND3X1_17 gnd vdd FILL
XFILL_9_NAND3X1_28 gnd vdd FILL
XFILL_9_NAND3X1_39 gnd vdd FILL
XFILL_15_BUFX4_19 gnd vdd FILL
XFILL_0_NOR3X1_5 gnd vdd FILL
XFILL_5_5_2 gnd vdd FILL
XFILL_4_0_1 gnd vdd FILL
XFILL_29_0_1 gnd vdd FILL
XFILL_2_NAND2X1_19 gnd vdd FILL
XFILL_33_DFFSR_5 gnd vdd FILL
XFILL_0_OAI21X1_4 gnd vdd FILL
XFILL_12_MUX2X1_150 gnd vdd FILL
XFILL_12_MUX2X1_161 gnd vdd FILL
XFILL_41_7_0 gnd vdd FILL
XFILL_12_MUX2X1_172 gnd vdd FILL
XFILL_13_4_2 gnd vdd FILL
XFILL_12_MUX2X1_183 gnd vdd FILL
XFILL_42_DFFSR_202 gnd vdd FILL
XFILL_12_MUX2X1_194 gnd vdd FILL
XFILL_42_DFFSR_213 gnd vdd FILL
XFILL_4_OAI21X1_3 gnd vdd FILL
XFILL_42_DFFSR_224 gnd vdd FILL
XFILL_42_DFFSR_235 gnd vdd FILL
XFILL_1_NOR2X1_50 gnd vdd FILL
XFILL_1_NOR2X1_61 gnd vdd FILL
XFILL_42_DFFSR_246 gnd vdd FILL
XFILL_42_DFFSR_257 gnd vdd FILL
XFILL_42_DFFSR_268 gnd vdd FILL
XFILL_1_NOR2X1_72 gnd vdd FILL
XFILL_1_NOR2X1_83 gnd vdd FILL
XFILL_1_NOR2X1_94 gnd vdd FILL
XFILL_46_DFFSR_201 gnd vdd FILL
XFILL_28_CLKBUF1_18 gnd vdd FILL
XFILL_46_DFFSR_212 gnd vdd FILL
XFILL_8_OAI21X1_2 gnd vdd FILL
XFILL_28_CLKBUF1_29 gnd vdd FILL
XFILL_46_DFFSR_223 gnd vdd FILL
XFILL_55_DFFSR_9 gnd vdd FILL
XFILL_46_DFFSR_234 gnd vdd FILL
XFILL_7_BUFX4_18 gnd vdd FILL
XFILL_5_NOR2X1_60 gnd vdd FILL
XFILL_7_BUFX4_29 gnd vdd FILL
XFILL_46_DFFSR_245 gnd vdd FILL
XFILL_5_NOR2X1_71 gnd vdd FILL
XFILL_46_DFFSR_256 gnd vdd FILL
XFILL_46_DFFSR_267 gnd vdd FILL
XFILL_5_NOR2X1_82 gnd vdd FILL
XFILL_73_DFFSR_101 gnd vdd FILL
XFILL_5_NOR2X1_93 gnd vdd FILL
XFILL_73_DFFSR_112 gnd vdd FILL
XFILL_6_AOI21X1_19 gnd vdd FILL
XFILL_73_DFFSR_123 gnd vdd FILL
XFILL_73_DFFSR_134 gnd vdd FILL
XFILL_73_DFFSR_145 gnd vdd FILL
XFILL_73_DFFSR_156 gnd vdd FILL
XFILL_9_NOR2X1_70 gnd vdd FILL
XFILL_73_DFFSR_167 gnd vdd FILL
XFILL_73_DFFSR_178 gnd vdd FILL
XFILL_9_NOR2X1_81 gnd vdd FILL
XFILL_9_NOR2X1_92 gnd vdd FILL
XFILL_77_DFFSR_100 gnd vdd FILL
XFILL_6_5 gnd vdd FILL
XFILL_73_DFFSR_189 gnd vdd FILL
XFILL_77_DFFSR_111 gnd vdd FILL
XFILL_9_NOR2X1_107 gnd vdd FILL
XFILL_77_DFFSR_122 gnd vdd FILL
XFILL_9_NOR2X1_118 gnd vdd FILL
XFILL_77_DFFSR_133 gnd vdd FILL
XFILL_77_DFFSR_144 gnd vdd FILL
XFILL_9_NOR2X1_129 gnd vdd FILL
XFILL_15_NAND3X1_20 gnd vdd FILL
XFILL_77_DFFSR_155 gnd vdd FILL
XFILL_15_NAND3X1_31 gnd vdd FILL
XFILL_77_DFFSR_166 gnd vdd FILL
XFILL_77_DFFSR_177 gnd vdd FILL
XFILL_15_NAND3X1_42 gnd vdd FILL
XFILL_15_NAND3X1_53 gnd vdd FILL
XFILL_77_DFFSR_188 gnd vdd FILL
XFILL_15_NAND3X1_64 gnd vdd FILL
XFILL_77_DFFSR_199 gnd vdd FILL
XFILL_15_NAND3X1_75 gnd vdd FILL
XFILL_35_CLKBUF1_20 gnd vdd FILL
XFILL_14_AND2X2_6 gnd vdd FILL
XFILL_15_NAND3X1_86 gnd vdd FILL
XFILL_35_CLKBUF1_31 gnd vdd FILL
XFILL_15_NAND3X1_97 gnd vdd FILL
XFILL_35_CLKBUF1_42 gnd vdd FILL
XFILL_63_3_2 gnd vdd FILL
XFILL_1_NAND2X1_5 gnd vdd FILL
XFILL_32_7_0 gnd vdd FILL
XFILL_11_BUFX4_12 gnd vdd FILL
XFILL_11_BUFX4_23 gnd vdd FILL
XFILL_11_BUFX4_34 gnd vdd FILL
XFILL_11_BUFX4_45 gnd vdd FILL
XFILL_5_NAND2X1_4 gnd vdd FILL
XFILL_11_BUFX4_56 gnd vdd FILL
XFILL_11_BUFX4_67 gnd vdd FILL
XFILL_11_BUFX4_78 gnd vdd FILL
XFILL_11_BUFX4_89 gnd vdd FILL
XFILL_6_OAI22X1_16 gnd vdd FILL
XFILL_6_OAI22X1_27 gnd vdd FILL
XFILL_14_NAND3X1_100 gnd vdd FILL
XFILL_1_MUX2X1_90 gnd vdd FILL
XFILL_14_NAND3X1_111 gnd vdd FILL
XFILL_6_OAI22X1_38 gnd vdd FILL
XFILL_14_NAND3X1_122 gnd vdd FILL
XDFFSR_15 DFFSR_15/Q DFFSR_88/CLK DFFSR_91/R vdd DFFSR_15/D gnd vdd DFFSR
XFILL_6_OAI22X1_49 gnd vdd FILL
XDFFSR_26 DFFSR_26/Q DFFSR_4/CLK DFFSR_26/R vdd DFFSR_26/D gnd vdd DFFSR
XFILL_9_NAND2X1_3 gnd vdd FILL
XFILL_13_DFFSR_201 gnd vdd FILL
XDFFSR_37 INVX1_21/A DFFSR_79/CLK DFFSR_48/R vdd MUX2X1_8/Y gnd vdd DFFSR
XFILL_13_DFFSR_212 gnd vdd FILL
XDFFSR_48 INVX1_15/A CLKBUF1_6/Y DFFSR_48/R vdd DFFSR_48/D gnd vdd DFFSR
XFILL_10_NAND3X1_1 gnd vdd FILL
XFILL_13_DFFSR_223 gnd vdd FILL
XDFFSR_59 DFFSR_59/Q DFFSR_97/CLK DFFSR_69/R vdd DFFSR_59/D gnd vdd DFFSR
XFILL_13_DFFSR_234 gnd vdd FILL
XFILL_13_DFFSR_245 gnd vdd FILL
XFILL_13_DFFSR_256 gnd vdd FILL
XFILL_13_DFFSR_267 gnd vdd FILL
XFILL_5_NAND3X1_70 gnd vdd FILL
XFILL_40_DFFSR_101 gnd vdd FILL
XFILL_5_NAND3X1_81 gnd vdd FILL
XFILL_5_NAND3X1_92 gnd vdd FILL
XFILL_17_DFFSR_200 gnd vdd FILL
XFILL_17_DFFSR_211 gnd vdd FILL
XFILL_9_NAND2X1_50 gnd vdd FILL
XFILL_40_DFFSR_112 gnd vdd FILL
XFILL_17_DFFSR_222 gnd vdd FILL
XFILL_9_NAND2X1_61 gnd vdd FILL
XFILL_40_DFFSR_123 gnd vdd FILL
XFILL_40_DFFSR_134 gnd vdd FILL
XFILL_5_INVX1_13 gnd vdd FILL
XFILL_9_NAND2X1_72 gnd vdd FILL
XFILL_17_DFFSR_233 gnd vdd FILL
XFILL_40_DFFSR_145 gnd vdd FILL
XFILL_9_NAND2X1_83 gnd vdd FILL
XFILL_22_10 gnd vdd FILL
XFILL_17_DFFSR_244 gnd vdd FILL
XCLKBUF1_13 BUFX4_10/Y gnd DFFSR_88/CLK vdd CLKBUF1
XFILL_5_INVX1_24 gnd vdd FILL
XFILL_5_NAND3X1_105 gnd vdd FILL
XFILL_40_DFFSR_156 gnd vdd FILL
XFILL_5_INVX1_35 gnd vdd FILL
XCLKBUF1_24 BUFX4_4/Y gnd CLKBUF1_24/Y vdd CLKBUF1
XFILL_17_DFFSR_255 gnd vdd FILL
XFILL_5_NAND3X1_116 gnd vdd FILL
XFILL_9_NAND2X1_94 gnd vdd FILL
XFILL_5_INVX1_46 gnd vdd FILL
XFILL_6_AND2X2_5 gnd vdd FILL
XFILL_40_DFFSR_167 gnd vdd FILL
XFILL_17_DFFSR_266 gnd vdd FILL
XFILL_40_DFFSR_178 gnd vdd FILL
XCLKBUF1_35 BUFX4_95/Y gnd DFFSR_52/CLK vdd CLKBUF1
XFILL_5_NAND3X1_127 gnd vdd FILL
XFILL_5_INVX1_57 gnd vdd FILL
XFILL_44_DFFSR_100 gnd vdd FILL
XFILL_40_DFFSR_189 gnd vdd FILL
XFILL_17_CLKBUF1_14 gnd vdd FILL
XFILL_5_INVX1_68 gnd vdd FILL
XFILL_44_DFFSR_111 gnd vdd FILL
XFILL_5_INVX1_79 gnd vdd FILL
XFILL_17_CLKBUF1_25 gnd vdd FILL
XFILL_44_DFFSR_122 gnd vdd FILL
XFILL_17_CLKBUF1_36 gnd vdd FILL
XFILL_5_AOI21X1_9 gnd vdd FILL
XFILL_44_DFFSR_133 gnd vdd FILL
XFILL_44_DFFSR_144 gnd vdd FILL
XFILL_12_AOI21X1_11 gnd vdd FILL
XFILL_44_DFFSR_155 gnd vdd FILL
XFILL_12_AOI21X1_22 gnd vdd FILL
XFILL_12_AOI21X1_33 gnd vdd FILL
XFILL_44_DFFSR_166 gnd vdd FILL
XFILL_12_AOI21X1_44 gnd vdd FILL
XFILL_2_DFFSR_4 gnd vdd FILL
XFILL_44_DFFSR_177 gnd vdd FILL
XFILL_44_DFFSR_188 gnd vdd FILL
XFILL_12_AOI21X1_55 gnd vdd FILL
XFILL_48_DFFSR_110 gnd vdd FILL
XFILL_44_DFFSR_199 gnd vdd FILL
XFILL_54_3_2 gnd vdd FILL
XFILL_12_AOI21X1_66 gnd vdd FILL
XFILL_15_DFFSR_2 gnd vdd FILL
XFILL_3_BUFX4_11 gnd vdd FILL
XFILL_12_AOI21X1_77 gnd vdd FILL
XFILL_48_DFFSR_121 gnd vdd FILL
XFILL_72_DFFSR_3 gnd vdd FILL
XFILL_48_DFFSR_132 gnd vdd FILL
XFILL_3_BUFX4_22 gnd vdd FILL
XFILL_9_AOI21X1_8 gnd vdd FILL
XFILL_48_DFFSR_143 gnd vdd FILL
XFILL_3_BUFX4_33 gnd vdd FILL
XFILL_48_DFFSR_154 gnd vdd FILL
XFILL_10_AOI22X1_6 gnd vdd FILL
XFILL_3_BUFX4_44 gnd vdd FILL
XFILL_48_DFFSR_165 gnd vdd FILL
XFILL_3_BUFX4_55 gnd vdd FILL
XFILL_48_DFFSR_176 gnd vdd FILL
XFILL_3_BUFX4_66 gnd vdd FILL
XFILL_48_DFFSR_187 gnd vdd FILL
XFILL_3_BUFX4_77 gnd vdd FILL
XFILL_48_DFFSR_198 gnd vdd FILL
XFILL_23_7_0 gnd vdd FILL
XFILL_3_BUFX4_88 gnd vdd FILL
XFILL_3_BUFX4_99 gnd vdd FILL
XFILL_10_BUFX2_8 gnd vdd FILL
XFILL_14_AOI22X1_5 gnd vdd FILL
XFILL_21_MUX2X1_9 gnd vdd FILL
XFILL_0_NAND3X1_101 gnd vdd FILL
XFILL_18_AOI22X1_4 gnd vdd FILL
XFILL_0_NAND3X1_112 gnd vdd FILL
XINVX1_109 DFFSR_57/Q gnd MUX2X1_96/A vdd INVX1
XFILL_37_DFFSR_6 gnd vdd FILL
XFILL_0_NAND3X1_123 gnd vdd FILL
XFILL_7_CLKBUF1_20 gnd vdd FILL
XFILL_29_DFFSR_13 gnd vdd FILL
XFILL_7_CLKBUF1_31 gnd vdd FILL
XFILL_29_DFFSR_24 gnd vdd FILL
XFILL_7_CLKBUF1_42 gnd vdd FILL
XFILL_15_MUX2X1_105 gnd vdd FILL
XFILL_29_DFFSR_35 gnd vdd FILL
XFILL_29_DFFSR_46 gnd vdd FILL
XFILL_15_MUX2X1_116 gnd vdd FILL
XFILL_29_DFFSR_57 gnd vdd FILL
XFILL_15_MUX2X1_127 gnd vdd FILL
XFILL_29_DFFSR_68 gnd vdd FILL
XFILL_15_MUX2X1_138 gnd vdd FILL
XFILL_15_MUX2X1_149 gnd vdd FILL
XFILL_2_AOI21X1_50 gnd vdd FILL
XFILL_29_DFFSR_79 gnd vdd FILL
XFILL_2_AOI21X1_61 gnd vdd FILL
XFILL_2_AOI21X1_72 gnd vdd FILL
XFILL_69_DFFSR_12 gnd vdd FILL
XFILL_12_OAI22X1_30 gnd vdd FILL
XFILL_12_OAI22X1_41 gnd vdd FILL
XFILL_69_DFFSR_23 gnd vdd FILL
XFILL_69_DFFSR_34 gnd vdd FILL
XFILL_69_DFFSR_45 gnd vdd FILL
XFILL_69_DFFSR_56 gnd vdd FILL
XFILL_69_DFFSR_67 gnd vdd FILL
XFILL_69_DFFSR_78 gnd vdd FILL
XFILL_5_NOR2X1_160 gnd vdd FILL
XFILL_69_DFFSR_89 gnd vdd FILL
XFILL_5_NOR2X1_171 gnd vdd FILL
XFILL_11_DFFSR_100 gnd vdd FILL
XFILL_5_NOR2X1_182 gnd vdd FILL
XFILL_5_NOR2X1_193 gnd vdd FILL
XFILL_11_DFFSR_111 gnd vdd FILL
XFILL_11_DFFSR_122 gnd vdd FILL
XFILL_11_DFFSR_133 gnd vdd FILL
XFILL_11_DFFSR_144 gnd vdd FILL
XFILL_38_DFFSR_11 gnd vdd FILL
XFILL_11_DFFSR_155 gnd vdd FILL
XFILL_38_DFFSR_22 gnd vdd FILL
XFILL_45_3_2 gnd vdd FILL
XFILL_38_DFFSR_33 gnd vdd FILL
XFILL_11_DFFSR_166 gnd vdd FILL
XFILL_0_CLKBUF1_9 gnd vdd FILL
XFILL_11_DFFSR_177 gnd vdd FILL
XFILL_38_DFFSR_44 gnd vdd FILL
XFILL_38_DFFSR_55 gnd vdd FILL
XFILL_11_DFFSR_188 gnd vdd FILL
XFILL_38_DFFSR_66 gnd vdd FILL
XFILL_15_DFFSR_110 gnd vdd FILL
XFILL_11_DFFSR_199 gnd vdd FILL
XFILL_38_DFFSR_77 gnd vdd FILL
XFILL_38_DFFSR_88 gnd vdd FILL
XFILL_15_DFFSR_121 gnd vdd FILL
XFILL_15_DFFSR_132 gnd vdd FILL
XFILL_15_DFFSR_143 gnd vdd FILL
XFILL_38_DFFSR_99 gnd vdd FILL
XFILL_78_DFFSR_10 gnd vdd FILL
XFILL_15_DFFSR_154 gnd vdd FILL
XFILL_78_DFFSR_21 gnd vdd FILL
XFILL_14_7_0 gnd vdd FILL
XFILL_22_MUX2X1_140 gnd vdd FILL
XFILL_78_DFFSR_32 gnd vdd FILL
XFILL_78_DFFSR_43 gnd vdd FILL
XFILL_15_DFFSR_165 gnd vdd FILL
XFILL_22_MUX2X1_151 gnd vdd FILL
XFILL_22_MUX2X1_162 gnd vdd FILL
XFILL_4_CLKBUF1_8 gnd vdd FILL
XFILL_15_DFFSR_176 gnd vdd FILL
XFILL_5_MUX2X1_100 gnd vdd FILL
XFILL_15_DFFSR_187 gnd vdd FILL
XFILL_78_DFFSR_54 gnd vdd FILL
XFILL_5_MUX2X1_111 gnd vdd FILL
XFILL_22_MUX2X1_173 gnd vdd FILL
XFILL_15_DFFSR_198 gnd vdd FILL
XFILL_78_DFFSR_65 gnd vdd FILL
XFILL_78_DFFSR_76 gnd vdd FILL
XFILL_5_MUX2X1_122 gnd vdd FILL
XFILL_19_DFFSR_120 gnd vdd FILL
XFILL_22_MUX2X1_184 gnd vdd FILL
XFILL_78_DFFSR_87 gnd vdd FILL
XFILL_5_MUX2X1_133 gnd vdd FILL
XFILL_19_DFFSR_131 gnd vdd FILL
XFILL_78_DFFSR_98 gnd vdd FILL
XFILL_5_MUX2X1_144 gnd vdd FILL
XFILL_19_DFFSR_142 gnd vdd FILL
XFILL_5_MUX2X1_155 gnd vdd FILL
XFILL_19_DFFSR_153 gnd vdd FILL
XFILL_0_BUFX4_103 gnd vdd FILL
XFILL_1_INVX1_50 gnd vdd FILL
XFILL_5_MUX2X1_166 gnd vdd FILL
XFILL_19_DFFSR_164 gnd vdd FILL
XFILL_1_INVX1_61 gnd vdd FILL
XFILL_5_MUX2X1_177 gnd vdd FILL
XFILL_8_CLKBUF1_7 gnd vdd FILL
XFILL_11_NOR3X1_11 gnd vdd FILL
XFILL_19_DFFSR_175 gnd vdd FILL
XFILL_1_INVX1_72 gnd vdd FILL
XFILL_1_INVX1_83 gnd vdd FILL
XFILL_19_DFFSR_186 gnd vdd FILL
XFILL_5_MUX2X1_188 gnd vdd FILL
XFILL_11_NOR3X1_22 gnd vdd FILL
XFILL_19_DFFSR_197 gnd vdd FILL
XFILL_11_NOR3X1_33 gnd vdd FILL
XFILL_47_DFFSR_20 gnd vdd FILL
XFILL_1_INVX1_94 gnd vdd FILL
XFILL_47_DFFSR_31 gnd vdd FILL
XFILL_61_DFFSR_200 gnd vdd FILL
XFILL_11_NOR3X1_44 gnd vdd FILL
XFILL_18_NOR3X1_6 gnd vdd FILL
XFILL_47_DFFSR_42 gnd vdd FILL
XFILL_61_DFFSR_211 gnd vdd FILL
XFILL_47_DFFSR_53 gnd vdd FILL
XFILL_61_DFFSR_222 gnd vdd FILL
XFILL_4_BUFX4_102 gnd vdd FILL
XFILL_47_DFFSR_64 gnd vdd FILL
XFILL_61_DFFSR_233 gnd vdd FILL
XFILL_47_DFFSR_75 gnd vdd FILL
XFILL_47_DFFSR_86 gnd vdd FILL
XFILL_61_DFFSR_244 gnd vdd FILL
XFILL_15_NOR3X1_10 gnd vdd FILL
XFILL_61_DFFSR_255 gnd vdd FILL
XFILL_47_DFFSR_97 gnd vdd FILL
XFILL_61_DFFSR_266 gnd vdd FILL
XFILL_15_NOR3X1_21 gnd vdd FILL
XFILL_15_NOR3X1_32 gnd vdd FILL
XFILL_87_DFFSR_30 gnd vdd FILL
XFILL_87_DFFSR_41 gnd vdd FILL
XFILL_15_NOR3X1_43 gnd vdd FILL
XFILL_65_DFFSR_210 gnd vdd FILL
XFILL_87_DFFSR_52 gnd vdd FILL
XFILL_87_DFFSR_63 gnd vdd FILL
XFILL_65_DFFSR_221 gnd vdd FILL
XFILL_8_BUFX4_101 gnd vdd FILL
XFILL_65_DFFSR_232 gnd vdd FILL
XFILL_87_DFFSR_74 gnd vdd FILL
XFILL_16_DFFSR_30 gnd vdd FILL
XFILL_65_DFFSR_243 gnd vdd FILL
XFILL_87_DFFSR_85 gnd vdd FILL
XFILL_16_DFFSR_41 gnd vdd FILL
XFILL_65_DFFSR_254 gnd vdd FILL
XFILL_87_DFFSR_96 gnd vdd FILL
XFILL_4_2 gnd vdd FILL
XFILL_16_DFFSR_52 gnd vdd FILL
XFILL_16_DFFSR_63 gnd vdd FILL
XFILL_65_DFFSR_265 gnd vdd FILL
XFILL_19_NOR3X1_20 gnd vdd FILL
XFILL_19_NOR3X1_31 gnd vdd FILL
XFILL_20_CLKBUF1_6 gnd vdd FILL
XFILL_16_DFFSR_74 gnd vdd FILL
XFILL_19_NOR3X1_42 gnd vdd FILL
XFILL_16_DFFSR_85 gnd vdd FILL
XFILL_60_4 gnd vdd FILL
XFILL_16_DFFSR_96 gnd vdd FILL
XFILL_69_DFFSR_220 gnd vdd FILL
XFILL_69_DFFSR_231 gnd vdd FILL
XFILL_56_DFFSR_40 gnd vdd FILL
XFILL_69_DFFSR_242 gnd vdd FILL
XFILL_27_NOR3X1_4 gnd vdd FILL
XFILL_56_DFFSR_51 gnd vdd FILL
XFILL_53_3 gnd vdd FILL
XFILL_69_DFFSR_253 gnd vdd FILL
XFILL_56_DFFSR_62 gnd vdd FILL
XFILL_69_DFFSR_264 gnd vdd FILL
XFILL_69_DFFSR_275 gnd vdd FILL
XFILL_56_DFFSR_73 gnd vdd FILL
XFILL_24_CLKBUF1_5 gnd vdd FILL
XFILL_64_6_0 gnd vdd FILL
XFILL_56_DFFSR_84 gnd vdd FILL
XFILL_36_3_2 gnd vdd FILL
XFILL_56_DFFSR_95 gnd vdd FILL
XFILL_46_2 gnd vdd FILL
XFILL_2_NOR2X1_15 gnd vdd FILL
XFILL_2_NOR2X1_26 gnd vdd FILL
XFILL_8_NAND3X1_14 gnd vdd FILL
XFILL_8_NAND3X1_25 gnd vdd FILL
XFILL_2_NOR2X1_37 gnd vdd FILL
XFILL_8_NAND3X1_36 gnd vdd FILL
XFILL_2_NOR2X1_48 gnd vdd FILL
XFILL_2_NOR2X1_59 gnd vdd FILL
XFILL_1_NOR2X1_5 gnd vdd FILL
XFILL_8_NAND3X1_47 gnd vdd FILL
XFILL_8_NAND3X1_58 gnd vdd FILL
XFILL_8_NAND3X1_69 gnd vdd FILL
XFILL_28_CLKBUF1_4 gnd vdd FILL
XFILL_6_NOR2X1_14 gnd vdd FILL
XFILL_25_DFFSR_50 gnd vdd FILL
XFILL_6_NOR2X1_25 gnd vdd FILL
XFILL_25_DFFSR_61 gnd vdd FILL
XFILL_6_NOR2X1_36 gnd vdd FILL
XFILL_25_DFFSR_72 gnd vdd FILL
XFILL_25_DFFSR_83 gnd vdd FILL
XFILL_6_NOR2X1_47 gnd vdd FILL
XFILL_6_NOR2X1_58 gnd vdd FILL
XFILL_10_OAI22X1_9 gnd vdd FILL
XFILL_6_NOR2X1_69 gnd vdd FILL
XFILL_25_DFFSR_94 gnd vdd FILL
XFILL_0_MUX2X1_3 gnd vdd FILL
XFILL_65_DFFSR_60 gnd vdd FILL
XFILL_65_DFFSR_71 gnd vdd FILL
XFILL_65_DFFSR_82 gnd vdd FILL
XFILL_14_OAI22X1_8 gnd vdd FILL
XFILL_65_DFFSR_93 gnd vdd FILL
XFILL_15_NAND3X1_101 gnd vdd FILL
XFILL_1_NAND2X1_16 gnd vdd FILL
XFILL_1_NAND2X1_27 gnd vdd FILL
XFILL_15_NAND3X1_112 gnd vdd FILL
XFILL_6_DFFSR_5 gnd vdd FILL
XFILL_15_NAND3X1_123 gnd vdd FILL
XFILL_1_NAND2X1_38 gnd vdd FILL
XFILL_19_DFFSR_3 gnd vdd FILL
XFILL_78_DFFSR_109 gnd vdd FILL
XFILL_1_NAND2X1_49 gnd vdd FILL
XFILL_76_DFFSR_4 gnd vdd FILL
XFILL_8_DFFSR_40 gnd vdd FILL
XFILL_8_DFFSR_51 gnd vdd FILL
XFILL_8_DFFSR_62 gnd vdd FILL
XFILL_18_OAI22X1_7 gnd vdd FILL
XFILL_8_DFFSR_73 gnd vdd FILL
XFILL_8_DFFSR_84 gnd vdd FILL
XFILL_8_DFFSR_95 gnd vdd FILL
XFILL_34_DFFSR_70 gnd vdd FILL
XFILL_34_DFFSR_81 gnd vdd FILL
XFILL_34_DFFSR_92 gnd vdd FILL
XFILL_11_MUX2X1_180 gnd vdd FILL
XFILL_11_MUX2X1_191 gnd vdd FILL
XFILL_32_DFFSR_210 gnd vdd FILL
XFILL_32_DFFSR_221 gnd vdd FILL
XFILL_32_DFFSR_232 gnd vdd FILL
XFILL_32_DFFSR_243 gnd vdd FILL
XFILL_6_NAND3X1_106 gnd vdd FILL
XFILL_32_DFFSR_254 gnd vdd FILL
XFILL_6_NAND3X1_117 gnd vdd FILL
XFILL_32_DFFSR_265 gnd vdd FILL
XFILL_74_DFFSR_80 gnd vdd FILL
XFILL_6_NAND3X1_128 gnd vdd FILL
XFILL_74_DFFSR_91 gnd vdd FILL
XFILL_27_CLKBUF1_15 gnd vdd FILL
XFILL_36_DFFSR_220 gnd vdd FILL
XFILL_27_CLKBUF1_26 gnd vdd FILL
XFILL_27_CLKBUF1_37 gnd vdd FILL
XFILL_36_DFFSR_231 gnd vdd FILL
XFILL_55_6_0 gnd vdd FILL
XFILL_36_DFFSR_242 gnd vdd FILL
XFILL_36_DFFSR_253 gnd vdd FILL
XFILL_2_3_2 gnd vdd FILL
XFILL_27_3_2 gnd vdd FILL
XFILL_36_DFFSR_264 gnd vdd FILL
XFILL_2_MUX2X1_11 gnd vdd FILL
XFILL_36_DFFSR_275 gnd vdd FILL
XFILL_2_MUX2X1_22 gnd vdd FILL
XFILL_2_MUX2X1_33 gnd vdd FILL
XFILL_2_MUX2X1_44 gnd vdd FILL
XFILL_5_AOI21X1_16 gnd vdd FILL
XFILL_63_DFFSR_120 gnd vdd FILL
XFILL_2_MUX2X1_55 gnd vdd FILL
XFILL_63_DFFSR_131 gnd vdd FILL
XFILL_2_MUX2X1_66 gnd vdd FILL
XFILL_5_AOI21X1_27 gnd vdd FILL
XFILL_43_DFFSR_90 gnd vdd FILL
XFILL_63_DFFSR_142 gnd vdd FILL
XFILL_2_MUX2X1_77 gnd vdd FILL
XFILL_63_DFFSR_153 gnd vdd FILL
XFILL_5_AOI21X1_38 gnd vdd FILL
XFILL_2_MUX2X1_88 gnd vdd FILL
XFILL_5_AOI21X1_49 gnd vdd FILL
XFILL_63_DFFSR_164 gnd vdd FILL
XFILL_2_MUX2X1_99 gnd vdd FILL
XFILL_6_MUX2X1_10 gnd vdd FILL
XFILL_6_MUX2X1_21 gnd vdd FILL
XFILL_63_DFFSR_175 gnd vdd FILL
XFILL_15_OAI22X1_18 gnd vdd FILL
XFILL_10_NAND3X1_130 gnd vdd FILL
XFILL_63_DFFSR_186 gnd vdd FILL
XFILL_15_OAI22X1_29 gnd vdd FILL
XFILL_63_DFFSR_197 gnd vdd FILL
XFILL_6_MUX2X1_32 gnd vdd FILL
XFILL_8_NOR2X1_104 gnd vdd FILL
XFILL_6_MUX2X1_43 gnd vdd FILL
XFILL_6_MUX2X1_54 gnd vdd FILL
XFILL_8_NOR2X1_115 gnd vdd FILL
XFILL_67_DFFSR_130 gnd vdd FILL
XFILL_6_MUX2X1_65 gnd vdd FILL
XFILL_8_NOR2X1_126 gnd vdd FILL
XFILL_67_DFFSR_141 gnd vdd FILL
XFILL_67_DFFSR_152 gnd vdd FILL
XFILL_6_MUX2X1_76 gnd vdd FILL
XFILL_8_NOR2X1_137 gnd vdd FILL
XFILL_0_BUFX4_5 gnd vdd FILL
XFILL_6_MUX2X1_87 gnd vdd FILL
XFILL_67_DFFSR_163 gnd vdd FILL
XFILL_10_2_2 gnd vdd FILL
XFILL_8_NOR2X1_148 gnd vdd FILL
XFILL_8_NOR2X1_159 gnd vdd FILL
XFILL_13_BUFX4_3 gnd vdd FILL
XFILL_6_MUX2X1_98 gnd vdd FILL
XFILL_67_DFFSR_174 gnd vdd FILL
XFILL_14_NAND3X1_50 gnd vdd FILL
XFILL_67_DFFSR_185 gnd vdd FILL
XFILL_14_NAND3X1_61 gnd vdd FILL
XFILL_67_DFFSR_196 gnd vdd FILL
XFILL_14_NAND3X1_72 gnd vdd FILL
XFILL_18_DFFSR_209 gnd vdd FILL
XFILL_14_NAND3X1_83 gnd vdd FILL
XFILL_15_NAND3X1_9 gnd vdd FILL
XFILL_14_NAND3X1_94 gnd vdd FILL
XFILL_1_NAND3X1_102 gnd vdd FILL
XFILL_1_NAND3X1_113 gnd vdd FILL
XFILL_1_NAND3X1_124 gnd vdd FILL
XFILL_45_DFFSR_109 gnd vdd FILL
XFILL_49_DFFSR_108 gnd vdd FILL
XFILL_49_DFFSR_119 gnd vdd FILL
XFILL_22_MUX2X1_30 gnd vdd FILL
XFILL_22_MUX2X1_41 gnd vdd FILL
XFILL_22_MUX2X1_52 gnd vdd FILL
XFILL_22_MUX2X1_63 gnd vdd FILL
XFILL_5_OAI22X1_13 gnd vdd FILL
XFILL_5_OAI22X1_24 gnd vdd FILL
XFILL_5_OAI22X1_35 gnd vdd FILL
XFILL_22_MUX2X1_74 gnd vdd FILL
XFILL_22_MUX2X1_85 gnd vdd FILL
XFILL_22_MUX2X1_96 gnd vdd FILL
XFILL_5_OAI22X1_46 gnd vdd FILL
XFILL_9_OAI21X1_15 gnd vdd FILL
XFILL_46_6_0 gnd vdd FILL
XFILL_9_OAI21X1_26 gnd vdd FILL
XFILL_18_3_2 gnd vdd FILL
XFILL_9_OAI21X1_37 gnd vdd FILL
XFILL_9_OAI21X1_48 gnd vdd FILL
XFILL_32_8 gnd vdd FILL
XFILL_60_1_2 gnd vdd FILL
XFILL_2_NOR2X1_204 gnd vdd FILL
XFILL_30_DFFSR_120 gnd vdd FILL
XFILL_30_DFFSR_131 gnd vdd FILL
XFILL_30_DFFSR_142 gnd vdd FILL
XFILL_8_NAND2X1_80 gnd vdd FILL
XFILL_30_DFFSR_153 gnd vdd FILL
XFILL_8_NAND2X1_91 gnd vdd FILL
XFILL_3_INVX8_3 gnd vdd FILL
XFILL_16_INVX8_1 gnd vdd FILL
XFILL_30_DFFSR_164 gnd vdd FILL
XFILL_30_DFFSR_175 gnd vdd FILL
XFILL_30_DFFSR_186 gnd vdd FILL
XFILL_16_CLKBUF1_11 gnd vdd FILL
XFILL_30_DFFSR_197 gnd vdd FILL
XFILL_16_CLKBUF1_22 gnd vdd FILL
XFILL_34_DFFSR_130 gnd vdd FILL
XFILL_16_CLKBUF1_33 gnd vdd FILL
XFILL_34_DFFSR_141 gnd vdd FILL
XFILL_34_DFFSR_152 gnd vdd FILL
XFILL_34_DFFSR_163 gnd vdd FILL
XFILL_11_AOI21X1_30 gnd vdd FILL
XFILL_34_DFFSR_174 gnd vdd FILL
XFILL_11_AOI21X1_41 gnd vdd FILL
XFILL_11_AOI21X1_52 gnd vdd FILL
XFILL_34_DFFSR_185 gnd vdd FILL
XFILL_20_DFFSR_3 gnd vdd FILL
XFILL_11_AOI21X1_63 gnd vdd FILL
XFILL_34_DFFSR_196 gnd vdd FILL
XFILL_11_AOI21X1_74 gnd vdd FILL
XFILL_38_DFFSR_140 gnd vdd FILL
XFILL_38_DFFSR_151 gnd vdd FILL
XFILL_58_DFFSR_1 gnd vdd FILL
XFILL_38_DFFSR_162 gnd vdd FILL
XFILL_38_DFFSR_173 gnd vdd FILL
XFILL_2_INVX1_17 gnd vdd FILL
XFILL_38_DFFSR_184 gnd vdd FILL
XFILL_2_INVX1_28 gnd vdd FILL
XFILL_30_NOR3X1_20 gnd vdd FILL
XFILL_30_NOR3X1_31 gnd vdd FILL
XFILL_38_DFFSR_195 gnd vdd FILL
XFILL_2_INVX1_39 gnd vdd FILL
XFILL_12_DFFSR_109 gnd vdd FILL
XFILL_30_NOR3X1_42 gnd vdd FILL
XFILL_80_DFFSR_220 gnd vdd FILL
XFILL_80_DFFSR_231 gnd vdd FILL
XFILL_80_DFFSR_242 gnd vdd FILL
XFILL_80_DFFSR_253 gnd vdd FILL
XFILL_80_DFFSR_264 gnd vdd FILL
XFILL_80_DFFSR_275 gnd vdd FILL
XFILL_16_DFFSR_108 gnd vdd FILL
XFILL_16_DFFSR_119 gnd vdd FILL
XFILL_84_DFFSR_230 gnd vdd FILL
XFILL_11_AOI21X1_4 gnd vdd FILL
XFILL_37_6_0 gnd vdd FILL
XFILL_0_BUFX4_15 gnd vdd FILL
XFILL_84_DFFSR_241 gnd vdd FILL
XFILL_0_BUFX4_26 gnd vdd FILL
XFILL_42_DFFSR_7 gnd vdd FILL
XFILL_0_BUFX4_37 gnd vdd FILL
XFILL_84_DFFSR_252 gnd vdd FILL
XFILL_0_BUFX4_48 gnd vdd FILL
XFILL_84_DFFSR_263 gnd vdd FILL
XFILL_84_DFFSR_274 gnd vdd FILL
XFILL_17_DFFSR_19 gnd vdd FILL
XFILL_0_BUFX4_59 gnd vdd FILL
XFILL_14_MUX2X1_102 gnd vdd FILL
XFILL_14_MUX2X1_113 gnd vdd FILL
XFILL_14_MUX2X1_124 gnd vdd FILL
XFILL_15_AOI21X1_3 gnd vdd FILL
XFILL_14_MUX2X1_135 gnd vdd FILL
XFILL_14_MUX2X1_146 gnd vdd FILL
XFILL_51_1_2 gnd vdd FILL
XFILL_0_INVX1_180 gnd vdd FILL
XFILL_14_MUX2X1_157 gnd vdd FILL
XFILL_14_MUX2X1_168 gnd vdd FILL
XFILL_0_INVX1_191 gnd vdd FILL
XFILL_1_AOI21X1_80 gnd vdd FILL
XFILL_57_DFFSR_18 gnd vdd FILL
XFILL_57_DFFSR_29 gnd vdd FILL
XFILL_14_MUX2X1_179 gnd vdd FILL
XFILL_62_DFFSR_209 gnd vdd FILL
XFILL_15_OAI21X1_40 gnd vdd FILL
XFILL_20_5_0 gnd vdd FILL
XFILL_4_INVX1_190 gnd vdd FILL
XFILL_16_NOR3X1_19 gnd vdd FILL
XFILL_4_NOR2X1_190 gnd vdd FILL
XFILL_66_DFFSR_208 gnd vdd FILL
XFILL_66_DFFSR_219 gnd vdd FILL
XFILL_26_DFFSR_17 gnd vdd FILL
XFILL_26_DFFSR_28 gnd vdd FILL
XFILL_26_DFFSR_39 gnd vdd FILL
XFILL_66_DFFSR_16 gnd vdd FILL
XFILL_66_DFFSR_27 gnd vdd FILL
XFILL_66_DFFSR_38 gnd vdd FILL
XFILL_66_DFFSR_49 gnd vdd FILL
XFILL_21_MUX2X1_170 gnd vdd FILL
XNAND3X1_15 DFFSR_40/Q BUFX4_5/Y NOR2X1_30/Y gnd NAND3X1_16/C vdd NAND3X1
XFILL_21_MUX2X1_181 gnd vdd FILL
XFILL_59_2_2 gnd vdd FILL
XNAND3X1_26 NOR3X1_44/Y NOR3X1_47/Y NOR3X1_43/Y gnd DFFSR_2/D vdd NAND3X1
XFILL_4_MUX2X1_130 gnd vdd FILL
XFILL_21_MUX2X1_192 gnd vdd FILL
XFILL_4_MUX2X1_141 gnd vdd FILL
XNAND3X1_37 OAI21X1_41/A INVX1_57/A NAND3X1_37/C gnd AOI22X1_3/D vdd NAND3X1
XNAND3X1_48 AOI22X1_1/A AOI22X1_1/B AND2X2_2/B gnd NOR3X1_49/B vdd NAND3X1
XFILL_9_DFFSR_18 gnd vdd FILL
XFILL_4_MUX2X1_152 gnd vdd FILL
XFILL_4_BUFX4_6 gnd vdd FILL
XFILL_4_MUX2X1_163 gnd vdd FILL
XNAND3X1_59 AND2X2_6/B AND2X2_6/A BUFX4_60/Y gnd OAI22X1_7/D vdd NAND3X1
XFILL_7_NAND3X1_107 gnd vdd FILL
XFILL_9_DFFSR_29 gnd vdd FILL
XFILL_4_MUX2X1_174 gnd vdd FILL
XFILL_4_MUX2X1_185 gnd vdd FILL
XFILL_7_NAND3X1_118 gnd vdd FILL
XFILL_35_DFFSR_15 gnd vdd FILL
XFILL_35_DFFSR_26 gnd vdd FILL
XFILL_35_DFFSR_37 gnd vdd FILL
XFILL_7_NAND3X1_129 gnd vdd FILL
XNOR2X1_15 NOR2X1_15/A NOR2X1_16/B gnd NOR2X1_15/Y vdd NOR2X1
XNOR2X1_26 NOR2X1_26/A NOR2X1_26/B gnd NOR2X1_26/Y vdd NOR2X1
XFILL_28_6_0 gnd vdd FILL
XNOR2X1_37 NOR3X1_51/C NOR2X1_37/B gnd NOR2X1_37/Y vdd NOR2X1
XFILL_3_6_0 gnd vdd FILL
XFILL_35_DFFSR_48 gnd vdd FILL
XFILL_35_DFFSR_59 gnd vdd FILL
XNOR2X1_48 NOR2X1_48/A NOR2X1_48/B gnd NOR2X1_48/Y vdd NOR2X1
XNOR2X1_59 OAI21X1_7/Y OAI21X1_6/Y gnd NOR2X1_59/Y vdd NOR2X1
XFILL_51_DFFSR_230 gnd vdd FILL
XFILL_51_DFFSR_241 gnd vdd FILL
XFILL_75_DFFSR_14 gnd vdd FILL
XFILL_51_DFFSR_252 gnd vdd FILL
XFILL_75_DFFSR_25 gnd vdd FILL
XFILL_51_DFFSR_263 gnd vdd FILL
XFILL_51_DFFSR_274 gnd vdd FILL
XFILL_75_DFFSR_36 gnd vdd FILL
XFILL_75_DFFSR_47 gnd vdd FILL
XFILL_18_MUX2X1_4 gnd vdd FILL
XFILL_42_1_2 gnd vdd FILL
XFILL_75_DFFSR_58 gnd vdd FILL
XFILL_75_DFFSR_69 gnd vdd FILL
XFILL_55_DFFSR_240 gnd vdd FILL
XFILL_55_DFFSR_251 gnd vdd FILL
XFILL_11_NAND3X1_120 gnd vdd FILL
XFILL_11_NAND3X1_131 gnd vdd FILL
XFILL_55_DFFSR_262 gnd vdd FILL
XFILL_10_CLKBUF1_3 gnd vdd FILL
XFILL_55_DFFSR_273 gnd vdd FILL
XFILL_10_NAND2X1_18 gnd vdd FILL
XFILL_11_5_0 gnd vdd FILL
XFILL_10_NAND2X1_29 gnd vdd FILL
XFILL_44_DFFSR_13 gnd vdd FILL
XFILL_9_BUFX4_70 gnd vdd FILL
XFILL_0_BUFX2_2 gnd vdd FILL
XFILL_44_DFFSR_24 gnd vdd FILL
XFILL_44_DFFSR_35 gnd vdd FILL
XFILL_9_BUFX4_81 gnd vdd FILL
XFILL_82_DFFSR_140 gnd vdd FILL
XFILL_9_BUFX4_92 gnd vdd FILL
XFILL_44_DFFSR_46 gnd vdd FILL
XFILL_44_DFFSR_57 gnd vdd FILL
XFILL_82_DFFSR_151 gnd vdd FILL
XFILL_82_DFFSR_162 gnd vdd FILL
XFILL_59_DFFSR_250 gnd vdd FILL
XFILL_44_DFFSR_68 gnd vdd FILL
XFILL_59_DFFSR_261 gnd vdd FILL
XFILL_59_DFFSR_272 gnd vdd FILL
XFILL_82_DFFSR_173 gnd vdd FILL
XFILL_44_DFFSR_79 gnd vdd FILL
XFILL_14_CLKBUF1_2 gnd vdd FILL
XFILL_82_DFFSR_184 gnd vdd FILL
XFILL_2_DFFSR_210 gnd vdd FILL
XFILL_84_DFFSR_12 gnd vdd FILL
XFILL_82_DFFSR_195 gnd vdd FILL
XFILL_33_DFFSR_208 gnd vdd FILL
XFILL_7_NAND3X1_11 gnd vdd FILL
XFILL_2_DFFSR_221 gnd vdd FILL
XFILL_33_DFFSR_219 gnd vdd FILL
XFILL_2_DFFSR_232 gnd vdd FILL
XFILL_84_DFFSR_23 gnd vdd FILL
XFILL_7_NAND3X1_22 gnd vdd FILL
XFILL_84_DFFSR_34 gnd vdd FILL
XFILL_2_DFFSR_243 gnd vdd FILL
XFILL_2_NAND3X1_103 gnd vdd FILL
XFILL_7_NAND3X1_33 gnd vdd FILL
XFILL_84_DFFSR_45 gnd vdd FILL
XFILL_84_DFFSR_56 gnd vdd FILL
XFILL_13_DFFSR_12 gnd vdd FILL
XFILL_2_DFFSR_254 gnd vdd FILL
XFILL_2_NAND3X1_114 gnd vdd FILL
XFILL_86_DFFSR_150 gnd vdd FILL
XFILL_7_NAND3X1_44 gnd vdd FILL
XFILL_86_DFFSR_161 gnd vdd FILL
XFILL_7_NAND3X1_55 gnd vdd FILL
XFILL_84_DFFSR_67 gnd vdd FILL
XFILL_2_DFFSR_265 gnd vdd FILL
XFILL_18_CLKBUF1_1 gnd vdd FILL
XFILL_86_DFFSR_172 gnd vdd FILL
XFILL_2_NAND3X1_125 gnd vdd FILL
XFILL_13_DFFSR_23 gnd vdd FILL
XFILL_7_NAND3X1_66 gnd vdd FILL
XFILL_84_DFFSR_78 gnd vdd FILL
XFILL_13_DFFSR_34 gnd vdd FILL
XFILL_84_DFFSR_89 gnd vdd FILL
XFILL_7_NAND3X1_77 gnd vdd FILL
XFILL_86_DFFSR_183 gnd vdd FILL
XFILL_13_DFFSR_45 gnd vdd FILL
XFILL_13_DFFSR_56 gnd vdd FILL
XFILL_60_DFFSR_108 gnd vdd FILL
XFILL_7_NAND3X1_88 gnd vdd FILL
XFILL_86_DFFSR_194 gnd vdd FILL
XFILL_37_DFFSR_207 gnd vdd FILL
XFILL_7_NAND3X1_99 gnd vdd FILL
XFILL_13_DFFSR_67 gnd vdd FILL
XFILL_6_DFFSR_220 gnd vdd FILL
XFILL_60_DFFSR_119 gnd vdd FILL
XFILL_37_DFFSR_218 gnd vdd FILL
XFILL_6_DFFSR_231 gnd vdd FILL
XFILL_13_DFFSR_78 gnd vdd FILL
XFILL_37_DFFSR_229 gnd vdd FILL
XFILL_13_DFFSR_89 gnd vdd FILL
XFILL_7_INVX8_4 gnd vdd FILL
XFILL_6_DFFSR_242 gnd vdd FILL
XFILL_53_DFFSR_11 gnd vdd FILL
XFILL_6_DFFSR_253 gnd vdd FILL
XFILL_53_DFFSR_22 gnd vdd FILL
XFILL_6_DFFSR_264 gnd vdd FILL
XFILL_6_DFFSR_275 gnd vdd FILL
XFILL_53_DFFSR_33 gnd vdd FILL
XFILL_24_NOR3X1_8 gnd vdd FILL
XFILL_53_DFFSR_44 gnd vdd FILL
XFILL_64_DFFSR_107 gnd vdd FILL
XFILL_53_DFFSR_55 gnd vdd FILL
XFILL_53_DFFSR_66 gnd vdd FILL
XFILL_53_DFFSR_77 gnd vdd FILL
XFILL_64_DFFSR_118 gnd vdd FILL
XFILL_64_DFFSR_129 gnd vdd FILL
XFILL_53_DFFSR_88 gnd vdd FILL
XFILL_53_DFFSR_99 gnd vdd FILL
XFILL_14_AOI21X1_18 gnd vdd FILL
XFILL_19_6_0 gnd vdd FILL
XMUX2X1_11 MUX2X1_8/A NOR3X1_4/A MUX2X1_14/S gnd DFFSR_32/D vdd MUX2X1
XFILL_0_NAND2X1_13 gnd vdd FILL
XMUX2X1_22 MUX2X1_6/B INVX1_36/Y MUX2X1_22/S gnd DFFSR_4/D vdd MUX2X1
XFILL_14_AOI21X1_29 gnd vdd FILL
XFILL_0_NAND2X1_24 gnd vdd FILL
XFILL_7_MUX2X1_19 gnd vdd FILL
XMUX2X1_33 MUX2X1_9/A INVX1_47/Y NOR2X1_20/Y gnd MUX2X1_33/Y vdd MUX2X1
XFILL_0_NAND2X1_35 gnd vdd FILL
XFILL_24_DFFSR_4 gnd vdd FILL
XNOR2X1_105 OAI21X1_29/Y OAI22X1_44/Y gnd NOR2X1_105/Y vdd NOR2X1
XFILL_68_DFFSR_106 gnd vdd FILL
XMUX2X1_44 INVX1_58/Y MUX2X1_7/B NAND2X1_6/Y gnd MUX2X1_44/Y vdd MUX2X1
XFILL_22_DFFSR_10 gnd vdd FILL
XFILL_0_NAND2X1_46 gnd vdd FILL
XFILL_81_DFFSR_5 gnd vdd FILL
XFILL_22_DFFSR_21 gnd vdd FILL
XFILL_0_NAND2X1_57 gnd vdd FILL
XFILL_68_DFFSR_117 gnd vdd FILL
XMUX2X1_55 INVX1_69/Y BUFX4_65/Y NAND2X1_9/Y gnd MUX2X1_55/Y vdd MUX2X1
XNOR2X1_116 BUFX2_8/A BUFX2_9/A gnd OAI21X1_37/B vdd NOR2X1
XMUX2X1_66 MUX2X1_66/A INVX1_80/Y NOR2X1_23/Y gnd MUX2X1_66/Y vdd MUX2X1
XNOR2X1_127 DFFSR_151/Q AOI21X1_3/B gnd AOI21X1_3/C vdd NOR2X1
XFILL_22_DFFSR_32 gnd vdd FILL
XFILL_0_NAND2X1_68 gnd vdd FILL
XMUX2X1_77 BUFX4_64/Y INVX1_91/Y NOR2X1_26/B gnd MUX2X1_77/Y vdd MUX2X1
XFILL_0_NAND2X1_79 gnd vdd FILL
XFILL_68_DFFSR_128 gnd vdd FILL
XNOR2X1_138 NOR2X1_138/A INVX1_218/Y gnd INVX1_8/A vdd NOR2X1
XMUX2X1_88 OAI22X1_7/A BUFX4_64/Y MUX2X1_91/S gnd MUX2X1_88/Y vdd MUX2X1
XFILL_22_DFFSR_43 gnd vdd FILL
XNOR2X1_149 DFFSR_98/Q NOR2X1_153/B gnd NOR2X1_149/Y vdd NOR2X1
XFILL_68_DFFSR_139 gnd vdd FILL
XFILL_11_OAI21X1_7 gnd vdd FILL
XFILL_0_INVX2_2 gnd vdd FILL
XFILL_22_DFFSR_54 gnd vdd FILL
XFILL_61_4_0 gnd vdd FILL
XMUX2X1_99 MUX2X1_99/A BUFX4_96/Y MUX2X1_99/S gnd DFFSR_90/D vdd MUX2X1
XFILL_22_DFFSR_65 gnd vdd FILL
XFILL_22_DFFSR_76 gnd vdd FILL
XFILL_33_1_2 gnd vdd FILL
XFILL_22_DFFSR_87 gnd vdd FILL
XFILL_23_4 gnd vdd FILL
XFILL_22_DFFSR_98 gnd vdd FILL
XFILL_7_NOR3X1_9 gnd vdd FILL
XFILL_62_DFFSR_20 gnd vdd FILL
XFILL_62_DFFSR_31 gnd vdd FILL
XFILL_62_DFFSR_42 gnd vdd FILL
XFILL_16_3 gnd vdd FILL
XFILL_3_AOI22X1_3 gnd vdd FILL
XFILL_15_OAI21X1_6 gnd vdd FILL
XFILL_62_DFFSR_53 gnd vdd FILL
XFILL_22_DFFSR_240 gnd vdd FILL
XFILL_62_DFFSR_64 gnd vdd FILL
XFILL_22_DFFSR_251 gnd vdd FILL
XFILL_62_DFFSR_75 gnd vdd FILL
XFILL_62_DFFSR_86 gnd vdd FILL
XFILL_22_DFFSR_262 gnd vdd FILL
XFILL_22_DFFSR_273 gnd vdd FILL
XFILL_62_DFFSR_97 gnd vdd FILL
XFILL_3_INVX1_202 gnd vdd FILL
XFILL_26_CLKBUF1_12 gnd vdd FILL
XFILL_3_INVX1_213 gnd vdd FILL
XDFFSR_3 DFFSR_3/Q DFFSR_5/CLK DFFSR_5/R vdd DFFSR_3/D gnd vdd DFFSR
XFILL_26_CLKBUF1_23 gnd vdd FILL
XFILL_5_DFFSR_11 gnd vdd FILL
XFILL_3_INVX1_224 gnd vdd FILL
XFILL_5_DFFSR_22 gnd vdd FILL
XFILL_26_CLKBUF1_34 gnd vdd FILL
XFILL_7_AOI22X1_2 gnd vdd FILL
XFILL_5_DFFSR_33 gnd vdd FILL
XFILL_46_DFFSR_8 gnd vdd FILL
XFILL_5_DFFSR_44 gnd vdd FILL
XFILL_5_DFFSR_55 gnd vdd FILL
XFILL_31_DFFSR_30 gnd vdd FILL
XFILL_26_DFFSR_250 gnd vdd FILL
XFILL_5_DFFSR_66 gnd vdd FILL
XFILL_0_AOI22X1_11 gnd vdd FILL
XFILL_31_DFFSR_41 gnd vdd FILL
XFILL_26_DFFSR_261 gnd vdd FILL
XFILL_5_DFFSR_77 gnd vdd FILL
XFILL_9_CLKBUF1_16 gnd vdd FILL
XFILL_26_DFFSR_272 gnd vdd FILL
XFILL_31_DFFSR_52 gnd vdd FILL
XFILL_5_DFFSR_88 gnd vdd FILL
XFILL_23_MUX2X1_17 gnd vdd FILL
XFILL_9_CLKBUF1_27 gnd vdd FILL
XFILL_7_INVX1_201 gnd vdd FILL
XFILL_31_DFFSR_63 gnd vdd FILL
XFILL_9_CLKBUF1_38 gnd vdd FILL
XFILL_7_INVX1_212 gnd vdd FILL
XFILL_5_DFFSR_99 gnd vdd FILL
XFILL_7_INVX1_223 gnd vdd FILL
XFILL_31_DFFSR_74 gnd vdd FILL
XFILL_23_MUX2X1_28 gnd vdd FILL
XFILL_4_AOI21X1_13 gnd vdd FILL
XFILL_31_DFFSR_85 gnd vdd FILL
XFILL_23_MUX2X1_39 gnd vdd FILL
XFILL_31_DFFSR_96 gnd vdd FILL
XFILL_4_AOI21X1_24 gnd vdd FILL
XFILL_4_AOI21X1_35 gnd vdd FILL
XFILL_53_DFFSR_150 gnd vdd FILL
XFILL_53_DFFSR_161 gnd vdd FILL
XFILL_4_AOI21X1_46 gnd vdd FILL
XFILL_71_DFFSR_40 gnd vdd FILL
XFILL_53_DFFSR_172 gnd vdd FILL
XFILL_14_OAI22X1_15 gnd vdd FILL
XFILL_4_AOI21X1_57 gnd vdd FILL
XFILL_71_DFFSR_51 gnd vdd FILL
XFILL_4_AOI21X1_68 gnd vdd FILL
XFILL_53_DFFSR_183 gnd vdd FILL
XFILL_71_DFFSR_62 gnd vdd FILL
XFILL_14_OAI22X1_26 gnd vdd FILL
XFILL_4_AOI21X1_79 gnd vdd FILL
XFILL_53_DFFSR_194 gnd vdd FILL
XFILL_14_OAI22X1_37 gnd vdd FILL
XFILL_71_DFFSR_73 gnd vdd FILL
XINVX1_18 INVX1_18/A gnd MUX2X1_5/A vdd INVX1
XFILL_7_NOR2X1_101 gnd vdd FILL
XFILL_14_OAI22X1_48 gnd vdd FILL
XFILL_71_DFFSR_84 gnd vdd FILL
XINVX1_29 INVX1_29/A gnd INVX1_29/Y vdd INVX1
XFILL_7_NOR2X1_112 gnd vdd FILL
XFILL_71_DFFSR_95 gnd vdd FILL
XFILL_7_NOR2X1_123 gnd vdd FILL
XFILL_7_NOR2X1_134 gnd vdd FILL
XFILL_57_DFFSR_160 gnd vdd FILL
XFILL_7_NOR2X1_145 gnd vdd FILL
XFILL_7_NOR2X1_156 gnd vdd FILL
XFILL_57_DFFSR_171 gnd vdd FILL
XFILL_7_NOR2X1_167 gnd vdd FILL
XFILL_7_NOR2X1_178 gnd vdd FILL
XFILL_57_DFFSR_182 gnd vdd FILL
XFILL_31_DFFSR_107 gnd vdd FILL
XFILL_57_DFFSR_193 gnd vdd FILL
XFILL_0_DFFSR_120 gnd vdd FILL
XFILL_11_NOR3X1_3 gnd vdd FILL
XFILL_7_NOR2X1_189 gnd vdd FILL
XNAND2X1_70 BUFX4_5/Y NOR2X1_29/Y gnd OAI22X1_26/D vdd NAND2X1
XFILL_0_DFFSR_131 gnd vdd FILL
XNAND2X1_81 NOR2X1_107/Y NOR2X1_106/Y gnd NOR3X1_47/B vdd NAND2X1
XFILL_31_DFFSR_118 gnd vdd FILL
XFILL_13_NAND3X1_80 gnd vdd FILL
XFILL_13_NAND3X1_91 gnd vdd FILL
XFILL_0_DFFSR_142 gnd vdd FILL
XFILL_31_DFFSR_129 gnd vdd FILL
XFILL_40_DFFSR_50 gnd vdd FILL
XFILL_0_DFFSR_153 gnd vdd FILL
XNAND2X1_92 INVX1_130/A INVX1_132/Y gnd NAND2X1_92/Y vdd NAND2X1
XFILL_40_DFFSR_61 gnd vdd FILL
XFILL_11_NOR2X1_206 gnd vdd FILL
XFILL_40_DFFSR_72 gnd vdd FILL
XFILL_0_DFFSR_164 gnd vdd FILL
XFILL_40_DFFSR_83 gnd vdd FILL
XFILL_0_DFFSR_175 gnd vdd FILL
XFILL_0_DFFSR_186 gnd vdd FILL
XFILL_40_DFFSR_94 gnd vdd FILL
XFILL_0_DFFSR_197 gnd vdd FILL
XFILL_35_DFFSR_106 gnd vdd FILL
XFILL_52_4_0 gnd vdd FILL
XFILL_35_DFFSR_117 gnd vdd FILL
XFILL_4_DFFSR_130 gnd vdd FILL
XFILL_24_1_2 gnd vdd FILL
XFILL_35_DFFSR_128 gnd vdd FILL
XFILL_4_DFFSR_141 gnd vdd FILL
XFILL_4_DFFSR_152 gnd vdd FILL
XFILL_80_DFFSR_60 gnd vdd FILL
XFILL_35_DFFSR_139 gnd vdd FILL
XFILL_4_DFFSR_163 gnd vdd FILL
XFILL_80_DFFSR_71 gnd vdd FILL
XFILL_80_DFFSR_82 gnd vdd FILL
XFILL_4_DFFSR_174 gnd vdd FILL
XFILL_80_DFFSR_93 gnd vdd FILL
XFILL_4_DFFSR_185 gnd vdd FILL
XFILL_4_DFFSR_196 gnd vdd FILL
XFILL_39_DFFSR_105 gnd vdd FILL
XFILL_7_MUX2X1_107 gnd vdd FILL
XFILL_7_MUX2X1_118 gnd vdd FILL
XFILL_39_DFFSR_116 gnd vdd FILL
XFILL_7_MUX2X1_129 gnd vdd FILL
XFILL_39_DFFSR_127 gnd vdd FILL
XFILL_8_DFFSR_140 gnd vdd FILL
XFILL_39_DFFSR_138 gnd vdd FILL
XFILL_8_DFFSR_151 gnd vdd FILL
XFILL_8_DFFSR_162 gnd vdd FILL
XFILL_39_DFFSR_149 gnd vdd FILL
XFILL_4_OAI22X1_10 gnd vdd FILL
XFILL_12_MUX2X1_60 gnd vdd FILL
XFILL_8_BUFX4_7 gnd vdd FILL
XFILL_12_MUX2X1_71 gnd vdd FILL
XFILL_8_DFFSR_173 gnd vdd FILL
XFILL_20_NOR3X1_1 gnd vdd FILL
XFILL_4_OAI22X1_21 gnd vdd FILL
XFILL_4_OAI22X1_32 gnd vdd FILL
XFILL_8_DFFSR_184 gnd vdd FILL
XFILL_12_MUX2X1_82 gnd vdd FILL
XFILL_0_NOR3X1_20 gnd vdd FILL
XFILL_4_OAI22X1_43 gnd vdd FILL
XFILL_12_MUX2X1_93 gnd vdd FILL
XFILL_31_NOR3X1_18 gnd vdd FILL
XFILL_0_NOR3X1_31 gnd vdd FILL
XFILL_8_DFFSR_195 gnd vdd FILL
XFILL_8_OAI21X1_12 gnd vdd FILL
XFILL_0_NOR3X1_42 gnd vdd FILL
XFILL_31_NOR3X1_29 gnd vdd FILL
XFILL_8_OAI21X1_23 gnd vdd FILL
XFILL_81_DFFSR_207 gnd vdd FILL
XFILL_8_OAI21X1_34 gnd vdd FILL
XFILL_81_DFFSR_218 gnd vdd FILL
XFILL_8_OAI21X1_45 gnd vdd FILL
XFILL_81_DFFSR_229 gnd vdd FILL
XFILL_16_MUX2X1_70 gnd vdd FILL
XFILL_16_MUX2X1_81 gnd vdd FILL
XFILL_16_MUX2X1_92 gnd vdd FILL
XFILL_4_NOR3X1_30 gnd vdd FILL
XFILL_4_NOR3X1_41 gnd vdd FILL
XFILL_4_NOR3X1_52 gnd vdd FILL
XFILL_85_DFFSR_206 gnd vdd FILL
XFILL_1_NOR2X1_201 gnd vdd FILL
XFILL_85_DFFSR_217 gnd vdd FILL
XFILL_85_DFFSR_228 gnd vdd FILL
XFILL_20_DFFSR_150 gnd vdd FILL
XFILL_85_DFFSR_239 gnd vdd FILL
XFILL_20_DFFSR_161 gnd vdd FILL
XFILL_3_NOR3X1_2 gnd vdd FILL
XFILL_20_DFFSR_172 gnd vdd FILL
XFILL_7_2_2 gnd vdd FILL
XFILL_1_INVX1_101 gnd vdd FILL
XFILL_1_INVX1_112 gnd vdd FILL
XFILL_20_DFFSR_183 gnd vdd FILL
XFILL_8_NOR3X1_40 gnd vdd FILL
XFILL_8_NOR3X1_51 gnd vdd FILL
XFILL_20_DFFSR_194 gnd vdd FILL
XFILL_1_INVX1_123 gnd vdd FILL
XFILL_15_CLKBUF1_30 gnd vdd FILL
XFILL_4_BUFX2_3 gnd vdd FILL
XFILL_1_INVX1_134 gnd vdd FILL
XFILL_1_INVX1_145 gnd vdd FILL
XFILL_15_CLKBUF1_41 gnd vdd FILL
XFILL_1_INVX1_156 gnd vdd FILL
XFILL_1_INVX1_167 gnd vdd FILL
XFILL_24_DFFSR_160 gnd vdd FILL
XFILL_8_NAND3X1_108 gnd vdd FILL
XFILL_24_DFFSR_171 gnd vdd FILL
XFILL_1_INVX1_178 gnd vdd FILL
XFILL_5_INVX1_100 gnd vdd FILL
XFILL_1_INVX1_189 gnd vdd FILL
XFILL_8_NAND3X1_119 gnd vdd FILL
XFILL_5_INVX1_111 gnd vdd FILL
XFILL_24_DFFSR_182 gnd vdd FILL
XFILL_5_INVX1_122 gnd vdd FILL
XFILL_24_DFFSR_193 gnd vdd FILL
XFILL_10_AOI21X1_60 gnd vdd FILL
XFILL_10_AOI21X1_71 gnd vdd FILL
XFILL_5_INVX1_133 gnd vdd FILL
XFILL_5_INVX1_144 gnd vdd FILL
XFILL_5_INVX1_155 gnd vdd FILL
XFILL_63_DFFSR_2 gnd vdd FILL
XFILL_5_INVX1_166 gnd vdd FILL
XFILL_43_4_0 gnd vdd FILL
XFILL_1_DFFSR_70 gnd vdd FILL
XFILL_28_DFFSR_170 gnd vdd FILL
XFILL_1_DFFSR_81 gnd vdd FILL
XFILL_5_INVX1_177 gnd vdd FILL
XFILL_5_INVX1_188 gnd vdd FILL
XFILL_1_DFFSR_92 gnd vdd FILL
XFILL_15_1_2 gnd vdd FILL
XFILL_28_DFFSR_181 gnd vdd FILL
XFILL_5_INVX1_199 gnd vdd FILL
XFILL_28_DFFSR_192 gnd vdd FILL
XFILL_20_NOR3X1_50 gnd vdd FILL
XFILL_12_NAND3X1_110 gnd vdd FILL
XFILL_12_NAND3X1_121 gnd vdd FILL
XFILL_70_DFFSR_250 gnd vdd FILL
XFILL_12_NAND3X1_132 gnd vdd FILL
XFILL_70_DFFSR_261 gnd vdd FILL
XFILL_70_DFFSR_272 gnd vdd FILL
XFILL_3_OAI22X1_6 gnd vdd FILL
XFILL_28_DFFSR_5 gnd vdd FILL
XFILL_74_DFFSR_260 gnd vdd FILL
XFILL_74_DFFSR_271 gnd vdd FILL
XFILL_85_DFFSR_6 gnd vdd FILL
XFILL_13_MUX2X1_110 gnd vdd FILL
XFILL_13_MUX2X1_121 gnd vdd FILL
XFILL_7_OAI22X1_5 gnd vdd FILL
XFILL_13_MUX2X1_132 gnd vdd FILL
XFILL_4_INVX2_3 gnd vdd FILL
XFILL_3_NAND3X1_104 gnd vdd FILL
XFILL_3_NAND3X1_115 gnd vdd FILL
XFILL_13_MUX2X1_143 gnd vdd FILL
XFILL_13_MUX2X1_154 gnd vdd FILL
XFILL_3_NAND3X1_126 gnd vdd FILL
XFILL_13_MUX2X1_165 gnd vdd FILL
XFILL_78_DFFSR_270 gnd vdd FILL
XFILL_13_MUX2X1_176 gnd vdd FILL
XFILL_13_MUX2X1_187 gnd vdd FILL
XFILL_52_DFFSR_206 gnd vdd FILL
XFILL_52_DFFSR_217 gnd vdd FILL
XFILL_52_DFFSR_228 gnd vdd FILL
XFILL_52_DFFSR_239 gnd vdd FILL
XFILL_2_INVX1_1 gnd vdd FILL
XFILL_56_DFFSR_205 gnd vdd FILL
XFILL_65_0_2 gnd vdd FILL
XFILL_56_DFFSR_216 gnd vdd FILL
XFILL_56_DFFSR_227 gnd vdd FILL
XFILL_56_DFFSR_238 gnd vdd FILL
XFILL_56_DFFSR_249 gnd vdd FILL
XFILL_83_DFFSR_105 gnd vdd FILL
XFILL_34_4_0 gnd vdd FILL
XFILL_83_DFFSR_116 gnd vdd FILL
XFILL_83_DFFSR_127 gnd vdd FILL
XFILL_83_DFFSR_138 gnd vdd FILL
XFILL_83_DFFSR_149 gnd vdd FILL
XFILL_21_1 gnd vdd FILL
XFILL_87_DFFSR_104 gnd vdd FILL
XFILL_3_DFFSR_208 gnd vdd FILL
XFILL_3_DFFSR_219 gnd vdd FILL
XFILL_87_DFFSR_115 gnd vdd FILL
XFILL_0_NAND3X1_8 gnd vdd FILL
XFILL_87_DFFSR_126 gnd vdd FILL
XFILL_87_DFFSR_137 gnd vdd FILL
XFILL_14_BUFX4_20 gnd vdd FILL
XFILL_14_BUFX4_31 gnd vdd FILL
XFILL_87_DFFSR_148 gnd vdd FILL
XFILL_3_MUX2X1_160 gnd vdd FILL
XFILL_14_BUFX4_42 gnd vdd FILL
XFILL_3_MUX2X1_171 gnd vdd FILL
XFILL_87_DFFSR_159 gnd vdd FILL
XFILL_14_BUFX4_53 gnd vdd FILL
XFILL_3_MUX2X1_182 gnd vdd FILL
XFILL_3_MUX2X1_193 gnd vdd FILL
XFILL_14_BUFX4_64 gnd vdd FILL
XDFFSR_210 BUFX2_7/A DFFSR_6/CLK DFFSR_6/R vdd NOR3X1_9/A gnd vdd DFFSR
XFILL_7_DFFSR_207 gnd vdd FILL
XFILL_4_NAND3X1_7 gnd vdd FILL
XDFFSR_221 BUFX2_8/A CLKBUF1_24/Y BUFX4_32/Y vdd INVX1_138/Y gnd vdd DFFSR
XFILL_14_BUFX4_75 gnd vdd FILL
XDFFSR_232 BUFX2_9/A CLKBUF1_24/Y BUFX4_32/Y vdd AND2X2_2/B gnd vdd DFFSR
XFILL_7_DFFSR_218 gnd vdd FILL
XFILL_14_BUFX4_86 gnd vdd FILL
XDFFSR_243 BUFX2_10/A DFFSR_84/CLK DFFSR_84/R vdd DFFSR_243/D gnd vdd DFFSR
XFILL_14_BUFX4_97 gnd vdd FILL
XFILL_7_DFFSR_229 gnd vdd FILL
XDFFSR_254 BUFX2_1/A DFFSR_93/CLK DFFSR_89/R vdd DFFSR_254/D gnd vdd DFFSR
XDFFSR_265 BUFX2_2/A DFFSR_70/CLK DFFSR_96/R vdd NAND3X1_4/Y gnd vdd DFFSR
XFILL_15_BUFX4_105 gnd vdd FILL
XFILL_41_DFFSR_260 gnd vdd FILL
XFILL_41_DFFSR_271 gnd vdd FILL
XFILL_8_NAND3X1_6 gnd vdd FILL
XFILL_45_DFFSR_270 gnd vdd FILL
XFILL_32_DFFSR_19 gnd vdd FILL
XFILL_9_AND2X2_2 gnd vdd FILL
XFILL_72_DFFSR_170 gnd vdd FILL
XFILL_56_0_2 gnd vdd FILL
XFILL_72_DFFSR_181 gnd vdd FILL
XFILL_72_DFFSR_18 gnd vdd FILL
XFILL_72_DFFSR_192 gnd vdd FILL
XFILL_23_DFFSR_205 gnd vdd FILL
XFILL_72_DFFSR_29 gnd vdd FILL
XFILL_23_DFFSR_216 gnd vdd FILL
XFILL_23_DFFSR_227 gnd vdd FILL
XFILL_15_MUX2X1_8 gnd vdd FILL
XFILL_6_NAND3X1_30 gnd vdd FILL
XFILL_23_DFFSR_238 gnd vdd FILL
XFILL_6_NAND3X1_41 gnd vdd FILL
XFILL_23_DFFSR_249 gnd vdd FILL
XFILL_25_4_0 gnd vdd FILL
XFILL_6_NAND3X1_52 gnd vdd FILL
XFILL_0_4_0 gnd vdd FILL
XFILL_6_NAND3X1_63 gnd vdd FILL
XFILL_76_DFFSR_180 gnd vdd FILL
XFILL_6_NAND3X1_74 gnd vdd FILL
XFILL_50_DFFSR_105 gnd vdd FILL
XFILL_6_NAND3X1_85 gnd vdd FILL
XFILL_76_DFFSR_191 gnd vdd FILL
XFILL_6_NAND3X1_96 gnd vdd FILL
XFILL_6_BUFX4_30 gnd vdd FILL
XFILL_27_DFFSR_204 gnd vdd FILL
XFILL_27_DFFSR_215 gnd vdd FILL
XFILL_6_BUFX4_41 gnd vdd FILL
XFILL_50_DFFSR_116 gnd vdd FILL
XFILL_6_BUFX4_52 gnd vdd FILL
XFILL_50_DFFSR_127 gnd vdd FILL
XFILL_27_DFFSR_226 gnd vdd FILL
XFILL_50_DFFSR_138 gnd vdd FILL
XFILL_6_BUFX4_63 gnd vdd FILL
XFILL_27_DFFSR_237 gnd vdd FILL
XFILL_50_DFFSR_149 gnd vdd FILL
XFILL_41_DFFSR_17 gnd vdd FILL
XFILL_6_BUFX4_74 gnd vdd FILL
XFILL_27_DFFSR_248 gnd vdd FILL
XFILL_41_DFFSR_28 gnd vdd FILL
XFILL_6_BUFX4_85 gnd vdd FILL
XFILL_41_DFFSR_39 gnd vdd FILL
XFILL_27_DFFSR_259 gnd vdd FILL
XFILL_6_BUFX4_96 gnd vdd FILL
XFILL_54_DFFSR_104 gnd vdd FILL
XFILL_8_BUFX2_4 gnd vdd FILL
XFILL_18_CLKBUF1_18 gnd vdd FILL
XFILL_54_DFFSR_115 gnd vdd FILL
XFILL_18_CLKBUF1_29 gnd vdd FILL
XFILL_54_DFFSR_126 gnd vdd FILL
XFILL_54_DFFSR_137 gnd vdd FILL
XFILL_81_DFFSR_16 gnd vdd FILL
XFILL_54_DFFSR_148 gnd vdd FILL
XFILL_13_AOI21X1_15 gnd vdd FILL
XFILL_81_DFFSR_27 gnd vdd FILL
XFILL_54_DFFSR_159 gnd vdd FILL
XFILL_81_DFFSR_38 gnd vdd FILL
XFILL_13_AOI21X1_26 gnd vdd FILL
XFILL_13_AOI21X1_37 gnd vdd FILL
XFILL_81_DFFSR_49 gnd vdd FILL
XFILL_10_DFFSR_16 gnd vdd FILL
XFILL_13_AOI21X1_48 gnd vdd FILL
XFILL_13_AOI21X1_59 gnd vdd FILL
XFILL_58_DFFSR_103 gnd vdd FILL
XFILL_58_DFFSR_114 gnd vdd FILL
XFILL_10_DFFSR_27 gnd vdd FILL
XFILL_10_DFFSR_38 gnd vdd FILL
XFILL_58_DFFSR_125 gnd vdd FILL
XFILL_10_DFFSR_49 gnd vdd FILL
XFILL_67_DFFSR_3 gnd vdd FILL
XFILL_58_DFFSR_136 gnd vdd FILL
XFILL_58_DFFSR_147 gnd vdd FILL
XFILL_58_DFFSR_158 gnd vdd FILL
XFILL_8_NOR2X1_9 gnd vdd FILL
XFILL_58_DFFSR_169 gnd vdd FILL
XFILL_1_DFFSR_107 gnd vdd FILL
XFILL_50_DFFSR_15 gnd vdd FILL
XFILL_50_DFFSR_26 gnd vdd FILL
XFILL_1_DFFSR_118 gnd vdd FILL
XFILL_50_DFFSR_37 gnd vdd FILL
XFILL_1_DFFSR_129 gnd vdd FILL
XFILL_8_5_0 gnd vdd FILL
XFILL_50_DFFSR_48 gnd vdd FILL
XFILL_50_DFFSR_59 gnd vdd FILL
XFILL_5_DFFSR_106 gnd vdd FILL
XFILL_12_DFFSR_270 gnd vdd FILL
XFILL_5_DFFSR_117 gnd vdd FILL
XFILL_7_MUX2X1_7 gnd vdd FILL
XFILL_25_CLKBUF1_20 gnd vdd FILL
XFILL_5_DFFSR_128 gnd vdd FILL
XFILL_25_CLKBUF1_31 gnd vdd FILL
XFILL_5_DFFSR_139 gnd vdd FILL
XFILL_47_0_2 gnd vdd FILL
XFILL_0_AOI21X1_2 gnd vdd FILL
XFILL_51_DFFSR_9 gnd vdd FILL
XFILL_25_CLKBUF1_42 gnd vdd FILL
XFILL_9_NAND3X1_109 gnd vdd FILL
XFILL_9_DFFSR_105 gnd vdd FILL
XFILL_8_CLKBUF1_13 gnd vdd FILL
XFILL_10_BUFX4_90 gnd vdd FILL
XFILL_8_CLKBUF1_24 gnd vdd FILL
XFILL_9_DFFSR_116 gnd vdd FILL
XFILL_13_MUX2X1_14 gnd vdd FILL
XFILL_13_MUX2X1_25 gnd vdd FILL
XFILL_9_DFFSR_127 gnd vdd FILL
XFILL_8_CLKBUF1_35 gnd vdd FILL
XFILL_16_4_0 gnd vdd FILL
XFILL_9_DFFSR_138 gnd vdd FILL
XFILL_16_MUX2X1_109 gnd vdd FILL
XFILL_3_AOI21X1_10 gnd vdd FILL
XFILL_13_MUX2X1_36 gnd vdd FILL
XFILL_9_DFFSR_149 gnd vdd FILL
XFILL_3_AOI21X1_21 gnd vdd FILL
XFILL_13_MUX2X1_47 gnd vdd FILL
XFILL_4_AOI21X1_1 gnd vdd FILL
XFILL_3_AOI21X1_32 gnd vdd FILL
XFILL_13_MUX2X1_58 gnd vdd FILL
XFILL_3_AOI21X1_43 gnd vdd FILL
XFILL_13_MUX2X1_69 gnd vdd FILL
XOAI21X1_13 INVX1_156/Y OAI21X1_3/B OAI21X1_13/C gnd NOR2X1_75/A vdd OAI21X1
XFILL_1_NOR3X1_18 gnd vdd FILL
XFILL_3_AOI21X1_54 gnd vdd FILL
XFILL_13_OAI22X1_12 gnd vdd FILL
XFILL_13_OAI22X1_23 gnd vdd FILL
XFILL_1_NOR3X1_29 gnd vdd FILL
XFILL_3_AOI21X1_65 gnd vdd FILL
XFILL_43_DFFSR_180 gnd vdd FILL
XOAI21X1_24 INVX1_209/Y OAI21X1_5/B OAI21X1_24/C gnd NOR2X1_94/A vdd OAI21X1
XFILL_17_MUX2X1_13 gnd vdd FILL
XFILL_3_AOI21X1_76 gnd vdd FILL
XFILL_13_OAI22X1_34 gnd vdd FILL
XOAI21X1_35 OAI21X1_35/A NOR2X1_20/A OAI21X1_48/A gnd OAI21X1_35/Y vdd OAI21X1
XFILL_43_DFFSR_191 gnd vdd FILL
XFILL_17_MUX2X1_24 gnd vdd FILL
XOAI21X1_46 NOR2X1_24/A OAI21X1_46/B OAI21X1_46/C gnd AOI22X1_3/B vdd OAI21X1
XFILL_13_OAI22X1_45 gnd vdd FILL
XFILL_17_MUX2X1_35 gnd vdd FILL
XFILL_6_NOR2X1_120 gnd vdd FILL
XFILL_17_MUX2X1_46 gnd vdd FILL
XFILL_17_MUX2X1_57 gnd vdd FILL
XFILL_6_NOR2X1_131 gnd vdd FILL
XFILL_17_MUX2X1_68 gnd vdd FILL
XFILL_2_DFFSR_15 gnd vdd FILL
XFILL_17_MUX2X1_79 gnd vdd FILL
XFILL_2_DFFSR_26 gnd vdd FILL
XFILL_13_NAND3X1_100 gnd vdd FILL
XFILL_6_NOR2X1_142 gnd vdd FILL
XFILL_6_NOR2X1_153 gnd vdd FILL
XFILL_2_DFFSR_37 gnd vdd FILL
XFILL_5_NOR3X1_17 gnd vdd FILL
XFILL_13_NAND3X1_111 gnd vdd FILL
XFILL_5_NOR3X1_28 gnd vdd FILL
XFILL_6_INVX1_2 gnd vdd FILL
XFILL_13_NAND3X1_122 gnd vdd FILL
XFILL_6_NOR2X1_164 gnd vdd FILL
XFILL_6_NOR2X1_175 gnd vdd FILL
XFILL_2_DFFSR_48 gnd vdd FILL
XFILL_5_NOR3X1_39 gnd vdd FILL
XFILL_21_DFFSR_104 gnd vdd FILL
XFILL_47_DFFSR_190 gnd vdd FILL
XFILL_2_DFFSR_59 gnd vdd FILL
XFILL_6_NOR2X1_186 gnd vdd FILL
XFILL_21_DFFSR_115 gnd vdd FILL
XFILL_6_NOR2X1_197 gnd vdd FILL
XFILL_21_DFFSR_126 gnd vdd FILL
XFILL_21_DFFSR_137 gnd vdd FILL
XFILL_21_DFFSR_148 gnd vdd FILL
XFILL_10_NOR2X1_203 gnd vdd FILL
XFILL_4_INVX1_80 gnd vdd FILL
XFILL_21_DFFSR_159 gnd vdd FILL
XFILL_4_INVX1_91 gnd vdd FILL
XFILL_9_NOR3X1_16 gnd vdd FILL
XFILL_9_NOR3X1_27 gnd vdd FILL
XFILL_9_NOR3X1_38 gnd vdd FILL
XFILL_9_NOR3X1_49 gnd vdd FILL
XFILL_25_DFFSR_103 gnd vdd FILL
XFILL_11_MUX2X1_1 gnd vdd FILL
XFILL_25_DFFSR_114 gnd vdd FILL
XFILL_23_MUX2X1_100 gnd vdd FILL
XFILL_25_DFFSR_125 gnd vdd FILL
XFILL_23_MUX2X1_111 gnd vdd FILL
XFILL_25_DFFSR_136 gnd vdd FILL
XFILL_23_MUX2X1_122 gnd vdd FILL
XFILL_25_DFFSR_147 gnd vdd FILL
XFILL_25_DFFSR_158 gnd vdd FILL
XFILL_23_MUX2X1_133 gnd vdd FILL
XFILL_4_NAND3X1_105 gnd vdd FILL
XFILL_23_MUX2X1_144 gnd vdd FILL
XFILL_4_NAND3X1_116 gnd vdd FILL
XFILL_25_DFFSR_169 gnd vdd FILL
XFILL_23_MUX2X1_155 gnd vdd FILL
XFILL_4_NAND3X1_127 gnd vdd FILL
XFILL_6_INVX1_109 gnd vdd FILL
XFILL_23_MUX2X1_166 gnd vdd FILL
XFILL_29_DFFSR_102 gnd vdd FILL
XFILL_6_MUX2X1_104 gnd vdd FILL
XFILL_23_MUX2X1_177 gnd vdd FILL
XFILL_6_MUX2X1_115 gnd vdd FILL
XFILL_29_DFFSR_113 gnd vdd FILL
XFILL_29_DFFSR_124 gnd vdd FILL
XFILL_23_MUX2X1_188 gnd vdd FILL
XFILL_6_MUX2X1_126 gnd vdd FILL
XFILL_6_MUX2X1_137 gnd vdd FILL
XFILL_29_DFFSR_135 gnd vdd FILL
XFILL_6_MUX2X1_148 gnd vdd FILL
XFILL_29_DFFSR_146 gnd vdd FILL
XFILL_29_DFFSR_157 gnd vdd FILL
XFILL_6_MUX2X1_159 gnd vdd FILL
XFILL_19_DFFSR_60 gnd vdd FILL
XFILL_29_DFFSR_168 gnd vdd FILL
XFILL_19_DFFSR_71 gnd vdd FILL
XFILL_66_3_0 gnd vdd FILL
XFILL_19_DFFSR_82 gnd vdd FILL
XFILL_29_DFFSR_179 gnd vdd FILL
XFILL_3_OAI22X1_40 gnd vdd FILL
XFILL_21_NOR3X1_15 gnd vdd FILL
XFILL_38_0_2 gnd vdd FILL
XFILL_3_OAI22X1_51 gnd vdd FILL
XFILL_19_DFFSR_93 gnd vdd FILL
XFILL_21_NOR3X1_26 gnd vdd FILL
XFILL_7_OAI21X1_20 gnd vdd FILL
XFILL_21_NOR3X1_37 gnd vdd FILL
XFILL_21_NOR3X1_48 gnd vdd FILL
XFILL_7_OAI21X1_31 gnd vdd FILL
XFILL_71_DFFSR_204 gnd vdd FILL
XFILL_71_DFFSR_215 gnd vdd FILL
XFILL_7_OAI21X1_42 gnd vdd FILL
XFILL_71_DFFSR_226 gnd vdd FILL
XFILL_71_DFFSR_237 gnd vdd FILL
XFILL_59_DFFSR_70 gnd vdd FILL
XFILL_71_DFFSR_248 gnd vdd FILL
XFILL_59_DFFSR_81 gnd vdd FILL
XFILL_25_NOR3X1_14 gnd vdd FILL
XFILL_59_DFFSR_92 gnd vdd FILL
XFILL_71_DFFSR_259 gnd vdd FILL
XFILL_25_NOR3X1_25 gnd vdd FILL
XFILL_25_NOR3X1_36 gnd vdd FILL
XFILL_25_NOR3X1_47 gnd vdd FILL
XFILL_4_NOR2X1_2 gnd vdd FILL
XFILL_75_DFFSR_203 gnd vdd FILL
XFILL_75_DFFSR_214 gnd vdd FILL
XFILL_50_7_1 gnd vdd FILL
XFILL_75_DFFSR_225 gnd vdd FILL
XFILL_75_DFFSR_236 gnd vdd FILL
XFILL_75_DFFSR_247 gnd vdd FILL
XFILL_29_NOR3X1_13 gnd vdd FILL
XFILL_75_DFFSR_258 gnd vdd FILL
XFILL_10_DFFSR_180 gnd vdd FILL
XFILL_75_DFFSR_269 gnd vdd FILL
XFILL_29_NOR3X1_24 gnd vdd FILL
XFILL_29_NOR3X1_35 gnd vdd FILL
XFILL_10_DFFSR_191 gnd vdd FILL
XFILL_79_DFFSR_202 gnd vdd FILL
XFILL_29_NOR3X1_46 gnd vdd FILL
XFILL_28_DFFSR_80 gnd vdd FILL
XFILL_79_DFFSR_213 gnd vdd FILL
XFILL_28_DFFSR_91 gnd vdd FILL
XFILL_79_DFFSR_224 gnd vdd FILL
XFILL_79_DFFSR_235 gnd vdd FILL
XFILL_79_DFFSR_246 gnd vdd FILL
XFILL_79_DFFSR_257 gnd vdd FILL
XFILL_79_DFFSR_268 gnd vdd FILL
XFILL_34_CLKBUF1_9 gnd vdd FILL
XFILL_14_DFFSR_190 gnd vdd FILL
XFILL_11_DFFSR_2 gnd vdd FILL
XFILL_68_DFFSR_90 gnd vdd FILL
XFILL_9_NAND3X1_18 gnd vdd FILL
XFILL_9_NAND3X1_29 gnd vdd FILL
XFILL_0_NOR3X1_6 gnd vdd FILL
XFILL_57_3_0 gnd vdd FILL
XFILL_29_0_2 gnd vdd FILL
XFILL_4_0_2 gnd vdd FILL
XFILL_33_DFFSR_6 gnd vdd FILL
XFILL_0_OAI21X1_5 gnd vdd FILL
XFILL_12_MUX2X1_140 gnd vdd FILL
XFILL_12_MUX2X1_151 gnd vdd FILL
XFILL_12_MUX2X1_162 gnd vdd FILL
XFILL_12_MUX2X1_173 gnd vdd FILL
XFILL_41_7_1 gnd vdd FILL
XFILL_12_MUX2X1_184 gnd vdd FILL
XFILL_40_2_0 gnd vdd FILL
XFILL_42_DFFSR_203 gnd vdd FILL
XFILL_42_DFFSR_214 gnd vdd FILL
XFILL_4_OAI21X1_4 gnd vdd FILL
XFILL_42_DFFSR_225 gnd vdd FILL
XFILL_42_DFFSR_236 gnd vdd FILL
XFILL_1_NOR2X1_40 gnd vdd FILL
XFILL_1_NOR2X1_51 gnd vdd FILL
XFILL_1_NOR2X1_62 gnd vdd FILL
XFILL_42_DFFSR_247 gnd vdd FILL
XFILL_42_DFFSR_258 gnd vdd FILL
XFILL_1_NOR2X1_73 gnd vdd FILL
XFILL_42_DFFSR_269 gnd vdd FILL
XFILL_1_NOR2X1_84 gnd vdd FILL
XFILL_1_NOR2X1_95 gnd vdd FILL
XFILL_46_DFFSR_202 gnd vdd FILL
XFILL_28_CLKBUF1_19 gnd vdd FILL
XFILL_46_DFFSR_213 gnd vdd FILL
XFILL_8_OAI21X1_3 gnd vdd FILL
XFILL_46_DFFSR_224 gnd vdd FILL
XFILL_46_DFFSR_235 gnd vdd FILL
XFILL_7_BUFX4_19 gnd vdd FILL
XFILL_46_DFFSR_246 gnd vdd FILL
XFILL_5_NOR2X1_50 gnd vdd FILL
XFILL_5_NOR2X1_61 gnd vdd FILL
XFILL_46_DFFSR_257 gnd vdd FILL
XFILL_5_NOR2X1_72 gnd vdd FILL
XFILL_46_DFFSR_268 gnd vdd FILL
XFILL_5_NOR2X1_83 gnd vdd FILL
XFILL_73_DFFSR_102 gnd vdd FILL
XFILL_5_NOR2X1_94 gnd vdd FILL
XFILL_73_DFFSR_113 gnd vdd FILL
XFILL_73_DFFSR_124 gnd vdd FILL
XFILL_73_DFFSR_135 gnd vdd FILL
XFILL_73_DFFSR_146 gnd vdd FILL
XFILL_73_DFFSR_157 gnd vdd FILL
XFILL_9_NOR2X1_60 gnd vdd FILL
XFILL_9_NOR2X1_71 gnd vdd FILL
XFILL_73_DFFSR_168 gnd vdd FILL
XFILL_73_DFFSR_179 gnd vdd FILL
XFILL_9_NOR2X1_82 gnd vdd FILL
XFILL_9_NOR2X1_93 gnd vdd FILL
XFILL_77_DFFSR_101 gnd vdd FILL
XFILL_6_6 gnd vdd FILL
XFILL_77_DFFSR_112 gnd vdd FILL
XFILL_9_NOR2X1_108 gnd vdd FILL
XFILL_77_DFFSR_123 gnd vdd FILL
XFILL_77_DFFSR_134 gnd vdd FILL
XFILL_9_NOR2X1_119 gnd vdd FILL
XFILL_77_DFFSR_145 gnd vdd FILL
XFILL_15_NAND3X1_10 gnd vdd FILL
XFILL_77_DFFSR_156 gnd vdd FILL
XFILL_15_NAND3X1_21 gnd vdd FILL
XFILL_48_3_0 gnd vdd FILL
XFILL_77_DFFSR_167 gnd vdd FILL
XFILL_15_NAND3X1_32 gnd vdd FILL
XFILL_77_DFFSR_178 gnd vdd FILL
XFILL_2_MUX2X1_190 gnd vdd FILL
XFILL_15_NAND3X1_43 gnd vdd FILL
XFILL_15_NAND3X1_54 gnd vdd FILL
XFILL_77_DFFSR_189 gnd vdd FILL
XFILL_15_NAND3X1_65 gnd vdd FILL
XFILL_35_CLKBUF1_10 gnd vdd FILL
XFILL_35_CLKBUF1_21 gnd vdd FILL
XFILL_15_NAND3X1_76 gnd vdd FILL
XFILL_14_AND2X2_7 gnd vdd FILL
XFILL_35_CLKBUF1_32 gnd vdd FILL
XFILL_15_NAND3X1_87 gnd vdd FILL
XFILL_15_NAND3X1_98 gnd vdd FILL
XFILL_1_NAND2X1_6 gnd vdd FILL
XFILL_32_7_1 gnd vdd FILL
XFILL_11_BUFX4_13 gnd vdd FILL
XFILL_11_BUFX4_24 gnd vdd FILL
XFILL_31_2_0 gnd vdd FILL
XFILL_11_BUFX4_35 gnd vdd FILL
XFILL_11_BUFX4_46 gnd vdd FILL
XFILL_5_NAND2X1_5 gnd vdd FILL
XFILL_11_BUFX4_57 gnd vdd FILL
XFILL_11_BUFX4_68 gnd vdd FILL
XFILL_11_BUFX4_79 gnd vdd FILL
XFILL_1_MUX2X1_80 gnd vdd FILL
XFILL_6_OAI22X1_17 gnd vdd FILL
XFILL_14_NAND3X1_101 gnd vdd FILL
XFILL_6_OAI22X1_28 gnd vdd FILL
XFILL_1_MUX2X1_91 gnd vdd FILL
XFILL_6_OAI22X1_39 gnd vdd FILL
XFILL_14_NAND3X1_112 gnd vdd FILL
XDFFSR_16 DFFSR_16/Q DFFSR_87/CLK DFFSR_87/R vdd DFFSR_16/D gnd vdd DFFSR
XFILL_14_NAND3X1_123 gnd vdd FILL
XFILL_9_NAND2X1_4 gnd vdd FILL
XDFFSR_27 INVX1_29/A CLKBUF1_6/Y DFFSR_48/R vdd DFFSR_27/D gnd vdd DFFSR
XFILL_13_DFFSR_202 gnd vdd FILL
XFILL_19_AOI22X1_10 gnd vdd FILL
XDFFSR_38 INVX1_22/A CLKBUF1_4/Y DFFSR_57/R vdd MUX2X1_9/Y gnd vdd DFFSR
XFILL_10_NAND3X1_2 gnd vdd FILL
XFILL_13_DFFSR_213 gnd vdd FILL
XDFFSR_49 INVX1_16/A DFFSR_79/CLK DFFSR_49/R vdd MUX2X1_3/Y gnd vdd DFFSR
XFILL_13_DFFSR_224 gnd vdd FILL
XFILL_13_DFFSR_235 gnd vdd FILL
XFILL_5_MUX2X1_90 gnd vdd FILL
XFILL_13_DFFSR_246 gnd vdd FILL
XFILL_5_NAND3X1_60 gnd vdd FILL
XFILL_13_DFFSR_257 gnd vdd FILL
XFILL_13_DFFSR_268 gnd vdd FILL
XFILL_5_NAND3X1_71 gnd vdd FILL
XFILL_40_DFFSR_102 gnd vdd FILL
XFILL_5_NAND3X1_82 gnd vdd FILL
XFILL_9_NAND2X1_40 gnd vdd FILL
XFILL_17_DFFSR_201 gnd vdd FILL
XFILL_5_NAND3X1_93 gnd vdd FILL
XFILL_9_NAND2X1_51 gnd vdd FILL
XFILL_14_NAND3X1_1 gnd vdd FILL
XFILL_40_DFFSR_113 gnd vdd FILL
XFILL_17_DFFSR_212 gnd vdd FILL
XFILL_40_DFFSR_124 gnd vdd FILL
XFILL_9_NAND2X1_62 gnd vdd FILL
XFILL_17_DFFSR_223 gnd vdd FILL
XFILL_17_DFFSR_234 gnd vdd FILL
XFILL_9_NAND2X1_73 gnd vdd FILL
XFILL_40_DFFSR_135 gnd vdd FILL
XFILL_5_INVX1_14 gnd vdd FILL
XFILL_40_DFFSR_146 gnd vdd FILL
XFILL_17_DFFSR_245 gnd vdd FILL
XFILL_9_NAND2X1_84 gnd vdd FILL
XFILL_5_INVX1_25 gnd vdd FILL
XFILL_22_11 gnd vdd FILL
XFILL_40_DFFSR_157 gnd vdd FILL
XFILL_5_INVX1_36 gnd vdd FILL
XCLKBUF1_14 BUFX4_95/Y gnd DFFSR_47/CLK vdd CLKBUF1
XFILL_9_NAND2X1_95 gnd vdd FILL
XFILL_5_NAND3X1_106 gnd vdd FILL
XCLKBUF1_25 BUFX4_84/Y gnd DFFSR_81/CLK vdd CLKBUF1
XFILL_5_NAND3X1_117 gnd vdd FILL
XFILL_40_DFFSR_168 gnd vdd FILL
XFILL_17_DFFSR_256 gnd vdd FILL
XCLKBUF1_36 BUFX4_10/Y gnd DFFSR_87/CLK vdd CLKBUF1
XFILL_5_NAND3X1_128 gnd vdd FILL
XFILL_17_DFFSR_267 gnd vdd FILL
XFILL_5_INVX1_47 gnd vdd FILL
XFILL_6_AND2X2_6 gnd vdd FILL
XFILL_40_DFFSR_179 gnd vdd FILL
XFILL_5_INVX1_58 gnd vdd FILL
XFILL_44_DFFSR_101 gnd vdd FILL
XFILL_5_INVX1_69 gnd vdd FILL
XFILL_17_CLKBUF1_15 gnd vdd FILL
XFILL_44_DFFSR_112 gnd vdd FILL
XFILL_17_CLKBUF1_26 gnd vdd FILL
XFILL_44_DFFSR_123 gnd vdd FILL
XFILL_39_3_0 gnd vdd FILL
XFILL_17_CLKBUF1_37 gnd vdd FILL
XFILL_44_DFFSR_134 gnd vdd FILL
XFILL_44_DFFSR_145 gnd vdd FILL
XFILL_12_AOI21X1_12 gnd vdd FILL
XFILL_44_DFFSR_156 gnd vdd FILL
XFILL_12_AOI21X1_23 gnd vdd FILL
XFILL_44_DFFSR_167 gnd vdd FILL
XFILL_12_AOI21X1_34 gnd vdd FILL
XFILL_44_DFFSR_178 gnd vdd FILL
XFILL_2_DFFSR_5 gnd vdd FILL
XFILL_12_AOI21X1_45 gnd vdd FILL
XBUFX4_90 BUFX4_92/A gnd BUFX4_90/Y vdd BUFX4
XFILL_48_DFFSR_100 gnd vdd FILL
XFILL_44_DFFSR_189 gnd vdd FILL
XFILL_12_AOI21X1_56 gnd vdd FILL
XFILL_15_DFFSR_3 gnd vdd FILL
XFILL_12_AOI21X1_67 gnd vdd FILL
XFILL_48_DFFSR_111 gnd vdd FILL
XFILL_3_BUFX4_12 gnd vdd FILL
XFILL_12_AOI21X1_78 gnd vdd FILL
XFILL_48_DFFSR_122 gnd vdd FILL
XFILL_72_DFFSR_4 gnd vdd FILL
XFILL_48_DFFSR_133 gnd vdd FILL
XFILL_3_BUFX4_23 gnd vdd FILL
XFILL_9_AOI21X1_9 gnd vdd FILL
XFILL_48_DFFSR_144 gnd vdd FILL
XFILL_3_BUFX4_34 gnd vdd FILL
XFILL_3_BUFX4_45 gnd vdd FILL
XFILL_48_DFFSR_155 gnd vdd FILL
XFILL_10_AOI22X1_7 gnd vdd FILL
XFILL_3_BUFX4_56 gnd vdd FILL
XFILL_48_DFFSR_166 gnd vdd FILL
XFILL_48_DFFSR_177 gnd vdd FILL
XFILL_3_BUFX4_67 gnd vdd FILL
XFILL_3_BUFX4_78 gnd vdd FILL
XFILL_48_DFFSR_188 gnd vdd FILL
XFILL_23_7_1 gnd vdd FILL
XFILL_48_DFFSR_199 gnd vdd FILL
XFILL_3_BUFX4_89 gnd vdd FILL
XFILL_22_2_0 gnd vdd FILL
XFILL_10_BUFX2_9 gnd vdd FILL
XFILL_14_AOI22X1_6 gnd vdd FILL
XFILL_0_NAND3X1_102 gnd vdd FILL
XFILL_0_NAND3X1_113 gnd vdd FILL
XFILL_18_AOI22X1_5 gnd vdd FILL
XFILL_0_NAND3X1_124 gnd vdd FILL
XFILL_37_DFFSR_7 gnd vdd FILL
XFILL_7_CLKBUF1_10 gnd vdd FILL
XFILL_7_CLKBUF1_21 gnd vdd FILL
XFILL_7_CLKBUF1_32 gnd vdd FILL
XFILL_29_DFFSR_14 gnd vdd FILL
XFILL_29_DFFSR_25 gnd vdd FILL
XFILL_29_DFFSR_36 gnd vdd FILL
XFILL_15_MUX2X1_106 gnd vdd FILL
XFILL_15_MUX2X1_117 gnd vdd FILL
XFILL_15_MUX2X1_128 gnd vdd FILL
XFILL_29_DFFSR_47 gnd vdd FILL
XFILL_29_DFFSR_58 gnd vdd FILL
XFILL_2_AOI21X1_40 gnd vdd FILL
XFILL_2_AOI21X1_51 gnd vdd FILL
XFILL_15_MUX2X1_139 gnd vdd FILL
XFILL_29_DFFSR_69 gnd vdd FILL
XFILL_12_OAI22X1_20 gnd vdd FILL
XFILL_2_AOI21X1_62 gnd vdd FILL
XFILL_12_OAI22X1_31 gnd vdd FILL
XFILL_2_AOI21X1_73 gnd vdd FILL
XFILL_69_DFFSR_13 gnd vdd FILL
XFILL_12_OAI22X1_42 gnd vdd FILL
XFILL_69_DFFSR_24 gnd vdd FILL
XFILL_69_DFFSR_35 gnd vdd FILL
XFILL_69_DFFSR_46 gnd vdd FILL
XFILL_69_DFFSR_57 gnd vdd FILL
XFILL_69_DFFSR_68 gnd vdd FILL
XFILL_5_NOR2X1_150 gnd vdd FILL
XFILL_69_DFFSR_79 gnd vdd FILL
XFILL_5_NOR2X1_161 gnd vdd FILL
XFILL_5_3_0 gnd vdd FILL
XFILL_5_NOR2X1_172 gnd vdd FILL
XFILL_11_DFFSR_101 gnd vdd FILL
XFILL_5_NOR2X1_183 gnd vdd FILL
XFILL_11_DFFSR_112 gnd vdd FILL
XFILL_5_NOR2X1_194 gnd vdd FILL
XFILL_11_DFFSR_123 gnd vdd FILL
XFILL_11_DFFSR_134 gnd vdd FILL
XFILL_38_DFFSR_12 gnd vdd FILL
XFILL_11_DFFSR_145 gnd vdd FILL
XFILL_11_DFFSR_156 gnd vdd FILL
XFILL_38_DFFSR_23 gnd vdd FILL
XFILL_11_DFFSR_167 gnd vdd FILL
XFILL_38_DFFSR_34 gnd vdd FILL
XFILL_38_DFFSR_45 gnd vdd FILL
XFILL_11_DFFSR_178 gnd vdd FILL
XFILL_38_DFFSR_56 gnd vdd FILL
XFILL_15_DFFSR_100 gnd vdd FILL
XFILL_11_DFFSR_189 gnd vdd FILL
XFILL_38_DFFSR_67 gnd vdd FILL
XFILL_15_DFFSR_111 gnd vdd FILL
XFILL_38_DFFSR_78 gnd vdd FILL
XFILL_15_DFFSR_122 gnd vdd FILL
XFILL_38_DFFSR_89 gnd vdd FILL
XFILL_15_DFFSR_133 gnd vdd FILL
XFILL_78_DFFSR_11 gnd vdd FILL
XFILL_15_DFFSR_144 gnd vdd FILL
XFILL_14_7_1 gnd vdd FILL
XFILL_22_MUX2X1_130 gnd vdd FILL
XFILL_15_DFFSR_155 gnd vdd FILL
XFILL_78_DFFSR_22 gnd vdd FILL
XFILL_22_MUX2X1_141 gnd vdd FILL
XFILL_15_DFFSR_166 gnd vdd FILL
XFILL_78_DFFSR_33 gnd vdd FILL
XFILL_15_DFFSR_177 gnd vdd FILL
XFILL_13_2_0 gnd vdd FILL
XFILL_22_MUX2X1_152 gnd vdd FILL
XFILL_78_DFFSR_44 gnd vdd FILL
XFILL_22_MUX2X1_163 gnd vdd FILL
XFILL_4_CLKBUF1_9 gnd vdd FILL
XFILL_78_DFFSR_55 gnd vdd FILL
XFILL_5_MUX2X1_101 gnd vdd FILL
XFILL_78_DFFSR_66 gnd vdd FILL
XFILL_15_DFFSR_188 gnd vdd FILL
XFILL_22_MUX2X1_174 gnd vdd FILL
XFILL_22_MUX2X1_185 gnd vdd FILL
XFILL_5_MUX2X1_112 gnd vdd FILL
XFILL_19_DFFSR_110 gnd vdd FILL
XFILL_15_DFFSR_199 gnd vdd FILL
XFILL_5_MUX2X1_123 gnd vdd FILL
XFILL_78_DFFSR_77 gnd vdd FILL
XFILL_19_DFFSR_121 gnd vdd FILL
XFILL_19_DFFSR_132 gnd vdd FILL
XFILL_78_DFFSR_88 gnd vdd FILL
XFILL_5_MUX2X1_134 gnd vdd FILL
XFILL_5_MUX2X1_145 gnd vdd FILL
XFILL_78_DFFSR_99 gnd vdd FILL
XFILL_19_DFFSR_143 gnd vdd FILL
XFILL_1_INVX1_40 gnd vdd FILL
XFILL_19_DFFSR_154 gnd vdd FILL
XFILL_5_MUX2X1_156 gnd vdd FILL
XFILL_0_BUFX4_104 gnd vdd FILL
XFILL_1_INVX1_51 gnd vdd FILL
XFILL_19_DFFSR_165 gnd vdd FILL
XFILL_5_MUX2X1_167 gnd vdd FILL
XFILL_8_CLKBUF1_8 gnd vdd FILL
XFILL_5_MUX2X1_178 gnd vdd FILL
XFILL_1_INVX1_62 gnd vdd FILL
XFILL_19_DFFSR_176 gnd vdd FILL
XFILL_5_MUX2X1_189 gnd vdd FILL
XFILL_19_DFFSR_187 gnd vdd FILL
XFILL_11_NOR3X1_12 gnd vdd FILL
XFILL_47_DFFSR_10 gnd vdd FILL
XFILL_1_INVX1_73 gnd vdd FILL
XFILL_47_DFFSR_21 gnd vdd FILL
XFILL_1_INVX1_84 gnd vdd FILL
XFILL_11_NOR3X1_23 gnd vdd FILL
XFILL_11_NOR3X1_34 gnd vdd FILL
XFILL_19_DFFSR_198 gnd vdd FILL
XFILL_1_INVX1_95 gnd vdd FILL
XFILL_47_DFFSR_32 gnd vdd FILL
XFILL_11_NOR3X1_45 gnd vdd FILL
XFILL_61_DFFSR_201 gnd vdd FILL
XFILL_47_DFFSR_43 gnd vdd FILL
XFILL_18_NOR3X1_7 gnd vdd FILL
XFILL_61_DFFSR_212 gnd vdd FILL
XFILL_47_DFFSR_54 gnd vdd FILL
XFILL_6_OAI21X1_50 gnd vdd FILL
XFILL_47_DFFSR_65 gnd vdd FILL
XFILL_61_DFFSR_223 gnd vdd FILL
XFILL_47_DFFSR_76 gnd vdd FILL
XFILL_61_DFFSR_234 gnd vdd FILL
XFILL_4_BUFX4_103 gnd vdd FILL
XFILL_61_DFFSR_245 gnd vdd FILL
XFILL_15_NOR3X1_11 gnd vdd FILL
XFILL_47_DFFSR_87 gnd vdd FILL
XFILL_47_DFFSR_98 gnd vdd FILL
XFILL_61_DFFSR_256 gnd vdd FILL
XFILL_61_DFFSR_267 gnd vdd FILL
XFILL_87_DFFSR_20 gnd vdd FILL
XFILL_15_NOR3X1_22 gnd vdd FILL
XFILL_15_NOR3X1_33 gnd vdd FILL
XFILL_87_DFFSR_31 gnd vdd FILL
XFILL_65_DFFSR_200 gnd vdd FILL
XFILL_15_NOR3X1_44 gnd vdd FILL
XFILL_87_DFFSR_42 gnd vdd FILL
XFILL_65_DFFSR_211 gnd vdd FILL
XFILL_87_DFFSR_53 gnd vdd FILL
XFILL_65_DFFSR_222 gnd vdd FILL
XFILL_16_DFFSR_20 gnd vdd FILL
XFILL_87_DFFSR_64 gnd vdd FILL
XFILL_65_DFFSR_233 gnd vdd FILL
XFILL_8_BUFX4_102 gnd vdd FILL
XFILL_16_DFFSR_31 gnd vdd FILL
XFILL_87_DFFSR_75 gnd vdd FILL
XFILL_87_DFFSR_86 gnd vdd FILL
XFILL_65_DFFSR_244 gnd vdd FILL
XFILL_19_NOR3X1_10 gnd vdd FILL
XFILL_4_3 gnd vdd FILL
XFILL_16_DFFSR_42 gnd vdd FILL
XFILL_65_DFFSR_255 gnd vdd FILL
XFILL_16_DFFSR_53 gnd vdd FILL
XFILL_87_DFFSR_97 gnd vdd FILL
XFILL_12_INVX8_1 gnd vdd FILL
XFILL_16_DFFSR_64 gnd vdd FILL
XFILL_65_DFFSR_266 gnd vdd FILL
XFILL_19_NOR3X1_21 gnd vdd FILL
XFILL_20_CLKBUF1_7 gnd vdd FILL
XFILL_16_DFFSR_75 gnd vdd FILL
XFILL_19_NOR3X1_32 gnd vdd FILL
XFILL_16_DFFSR_86 gnd vdd FILL
XFILL_19_NOR3X1_43 gnd vdd FILL
XFILL_69_DFFSR_210 gnd vdd FILL
XFILL_60_5 gnd vdd FILL
XFILL_16_DFFSR_97 gnd vdd FILL
XFILL_69_DFFSR_221 gnd vdd FILL
XFILL_56_DFFSR_30 gnd vdd FILL
XFILL_69_DFFSR_232 gnd vdd FILL
XFILL_69_DFFSR_243 gnd vdd FILL
XFILL_56_DFFSR_41 gnd vdd FILL
XFILL_27_NOR3X1_5 gnd vdd FILL
XFILL_69_DFFSR_254 gnd vdd FILL
XFILL_53_4 gnd vdd FILL
XFILL_56_DFFSR_52 gnd vdd FILL
XFILL_56_DFFSR_63 gnd vdd FILL
XFILL_69_DFFSR_265 gnd vdd FILL
XFILL_24_CLKBUF1_6 gnd vdd FILL
XFILL_56_DFFSR_74 gnd vdd FILL
XFILL_64_6_1 gnd vdd FILL
XFILL_56_DFFSR_85 gnd vdd FILL
XFILL_46_3 gnd vdd FILL
XFILL_56_DFFSR_96 gnd vdd FILL
XFILL_2_NOR2X1_16 gnd vdd FILL
XFILL_63_1_0 gnd vdd FILL
XFILL_8_NAND3X1_15 gnd vdd FILL
XFILL_2_NOR2X1_27 gnd vdd FILL
XFILL_8_NAND3X1_26 gnd vdd FILL
XFILL_2_NOR2X1_38 gnd vdd FILL
XFILL_1_NOR2X1_6 gnd vdd FILL
XFILL_8_NAND3X1_37 gnd vdd FILL
XFILL_2_NOR2X1_49 gnd vdd FILL
XFILL_8_NAND3X1_48 gnd vdd FILL
XFILL_54_DFFSR_1 gnd vdd FILL
XFILL_8_NAND3X1_59 gnd vdd FILL
XFILL_28_CLKBUF1_5 gnd vdd FILL
XFILL_25_DFFSR_40 gnd vdd FILL
XFILL_25_DFFSR_51 gnd vdd FILL
XFILL_6_NOR2X1_15 gnd vdd FILL
XFILL_6_NOR2X1_26 gnd vdd FILL
XFILL_6_NOR2X1_37 gnd vdd FILL
XFILL_25_DFFSR_62 gnd vdd FILL
XFILL_25_DFFSR_73 gnd vdd FILL
XFILL_25_DFFSR_84 gnd vdd FILL
XFILL_6_NOR2X1_48 gnd vdd FILL
XFILL_25_DFFSR_95 gnd vdd FILL
XFILL_6_NOR2X1_59 gnd vdd FILL
XFILL_0_MUX2X1_4 gnd vdd FILL
XFILL_65_DFFSR_50 gnd vdd FILL
XFILL_65_DFFSR_61 gnd vdd FILL
XFILL_65_DFFSR_72 gnd vdd FILL
XFILL_65_DFFSR_83 gnd vdd FILL
XFILL_15_NAND3X1_102 gnd vdd FILL
XFILL_65_DFFSR_94 gnd vdd FILL
XFILL_14_OAI22X1_9 gnd vdd FILL
XFILL_1_NAND2X1_17 gnd vdd FILL
XFILL_15_NAND3X1_113 gnd vdd FILL
XFILL_1_NAND2X1_28 gnd vdd FILL
XFILL_6_DFFSR_6 gnd vdd FILL
XFILL_15_NAND3X1_124 gnd vdd FILL
XFILL_1_NAND2X1_39 gnd vdd FILL
XFILL_19_DFFSR_4 gnd vdd FILL
XFILL_8_DFFSR_30 gnd vdd FILL
XFILL_8_DFFSR_41 gnd vdd FILL
XFILL_76_DFFSR_5 gnd vdd FILL
XFILL_8_DFFSR_52 gnd vdd FILL
XFILL_8_DFFSR_63 gnd vdd FILL
XFILL_18_OAI22X1_8 gnd vdd FILL
XFILL_8_DFFSR_74 gnd vdd FILL
XFILL_8_DFFSR_85 gnd vdd FILL
XFILL_34_DFFSR_60 gnd vdd FILL
XFILL_8_DFFSR_96 gnd vdd FILL
XFILL_34_DFFSR_71 gnd vdd FILL
XFILL_11_MUX2X1_170 gnd vdd FILL
XFILL_34_DFFSR_82 gnd vdd FILL
XFILL_11_MUX2X1_181 gnd vdd FILL
XFILL_34_DFFSR_93 gnd vdd FILL
XFILL_32_DFFSR_200 gnd vdd FILL
XFILL_11_MUX2X1_192 gnd vdd FILL
XFILL_32_DFFSR_211 gnd vdd FILL
XFILL_32_DFFSR_222 gnd vdd FILL
XFILL_32_DFFSR_233 gnd vdd FILL
XFILL_32_DFFSR_244 gnd vdd FILL
XFILL_6_NAND3X1_107 gnd vdd FILL
XFILL_32_DFFSR_255 gnd vdd FILL
XFILL_6_NAND3X1_118 gnd vdd FILL
XFILL_74_DFFSR_70 gnd vdd FILL
XFILL_6_NAND3X1_129 gnd vdd FILL
XFILL_74_DFFSR_81 gnd vdd FILL
XFILL_32_DFFSR_266 gnd vdd FILL
XFILL_74_DFFSR_92 gnd vdd FILL
XFILL_27_CLKBUF1_16 gnd vdd FILL
XFILL_36_DFFSR_210 gnd vdd FILL
XFILL_27_CLKBUF1_27 gnd vdd FILL
XFILL_27_CLKBUF1_38 gnd vdd FILL
XFILL_36_DFFSR_221 gnd vdd FILL
XFILL_36_DFFSR_232 gnd vdd FILL
XFILL_36_DFFSR_243 gnd vdd FILL
XFILL_55_6_1 gnd vdd FILL
XFILL_36_DFFSR_254 gnd vdd FILL
XFILL_54_1_0 gnd vdd FILL
XFILL_2_MUX2X1_12 gnd vdd FILL
XFILL_36_DFFSR_265 gnd vdd FILL
XFILL_2_MUX2X1_23 gnd vdd FILL
XFILL_2_MUX2X1_34 gnd vdd FILL
XFILL_63_DFFSR_110 gnd vdd FILL
XFILL_2_MUX2X1_45 gnd vdd FILL
XFILL_63_DFFSR_121 gnd vdd FILL
XFILL_43_DFFSR_80 gnd vdd FILL
XFILL_63_DFFSR_132 gnd vdd FILL
XFILL_5_AOI21X1_17 gnd vdd FILL
XFILL_2_MUX2X1_56 gnd vdd FILL
XFILL_43_DFFSR_91 gnd vdd FILL
XFILL_5_AOI21X1_28 gnd vdd FILL
XFILL_2_MUX2X1_67 gnd vdd FILL
XFILL_63_DFFSR_143 gnd vdd FILL
XFILL_2_MUX2X1_78 gnd vdd FILL
XFILL_5_AOI21X1_39 gnd vdd FILL
XFILL_63_DFFSR_154 gnd vdd FILL
XFILL_63_DFFSR_165 gnd vdd FILL
XFILL_10_NAND3X1_120 gnd vdd FILL
XFILL_2_MUX2X1_89 gnd vdd FILL
XFILL_10_NAND3X1_131 gnd vdd FILL
XFILL_15_OAI22X1_19 gnd vdd FILL
XFILL_6_MUX2X1_11 gnd vdd FILL
XFILL_63_DFFSR_176 gnd vdd FILL
XFILL_6_MUX2X1_22 gnd vdd FILL
XFILL_63_DFFSR_187 gnd vdd FILL
XFILL_6_MUX2X1_33 gnd vdd FILL
XFILL_63_DFFSR_198 gnd vdd FILL
XFILL_6_MUX2X1_44 gnd vdd FILL
XFILL_8_NOR2X1_105 gnd vdd FILL
XFILL_67_DFFSR_120 gnd vdd FILL
XFILL_67_DFFSR_131 gnd vdd FILL
XFILL_6_MUX2X1_55 gnd vdd FILL
XFILL_8_NOR2X1_116 gnd vdd FILL
XFILL_83_DFFSR_90 gnd vdd FILL
XFILL_67_DFFSR_142 gnd vdd FILL
XFILL_6_MUX2X1_66 gnd vdd FILL
XFILL_8_NOR2X1_127 gnd vdd FILL
XFILL_6_MUX2X1_77 gnd vdd FILL
XFILL_8_NOR2X1_138 gnd vdd FILL
XFILL_6_MUX2X1_88 gnd vdd FILL
XFILL_67_DFFSR_153 gnd vdd FILL
XFILL_0_BUFX4_6 gnd vdd FILL
XFILL_8_NOR2X1_149 gnd vdd FILL
XFILL_67_DFFSR_164 gnd vdd FILL
XFILL_13_BUFX4_4 gnd vdd FILL
XFILL_6_MUX2X1_99 gnd vdd FILL
XFILL_67_DFFSR_175 gnd vdd FILL
XFILL_14_NAND3X1_40 gnd vdd FILL
XFILL_12_DFFSR_90 gnd vdd FILL
XFILL_67_DFFSR_186 gnd vdd FILL
XFILL_14_NAND3X1_51 gnd vdd FILL
XFILL_14_NAND3X1_62 gnd vdd FILL
XFILL_67_DFFSR_197 gnd vdd FILL
XFILL_14_NAND3X1_73 gnd vdd FILL
XFILL_14_NAND3X1_84 gnd vdd FILL
XFILL_14_NAND3X1_95 gnd vdd FILL
XFILL_34_CLKBUF1_40 gnd vdd FILL
XFILL_1_NAND3X1_103 gnd vdd FILL
XFILL_1_NAND3X1_114 gnd vdd FILL
XFILL_1_NAND3X1_125 gnd vdd FILL
XFILL_49_DFFSR_109 gnd vdd FILL
XFILL_22_MUX2X1_20 gnd vdd FILL
XFILL_22_MUX2X1_31 gnd vdd FILL
XFILL_22_MUX2X1_42 gnd vdd FILL
XFILL_22_MUX2X1_53 gnd vdd FILL
XFILL_22_MUX2X1_64 gnd vdd FILL
XFILL_5_OAI22X1_14 gnd vdd FILL
XFILL_22_MUX2X1_75 gnd vdd FILL
XFILL_5_OAI22X1_25 gnd vdd FILL
XFILL_22_MUX2X1_86 gnd vdd FILL
XFILL_5_OAI22X1_36 gnd vdd FILL
XFILL_5_OAI22X1_47 gnd vdd FILL
XFILL_22_MUX2X1_97 gnd vdd FILL
XFILL_46_6_1 gnd vdd FILL
XFILL_9_OAI21X1_16 gnd vdd FILL
XFILL_9_OAI21X1_27 gnd vdd FILL
XFILL_45_1_0 gnd vdd FILL
XFILL_9_OAI21X1_38 gnd vdd FILL
XFILL_9_OAI21X1_49 gnd vdd FILL
XFILL_32_9 gnd vdd FILL
XFILL_30_DFFSR_110 gnd vdd FILL
XFILL_4_NAND3X1_90 gnd vdd FILL
XFILL_2_NOR2X1_205 gnd vdd FILL
XFILL_30_DFFSR_121 gnd vdd FILL
XFILL_30_DFFSR_132 gnd vdd FILL
XFILL_8_NAND2X1_70 gnd vdd FILL
XFILL_30_DFFSR_143 gnd vdd FILL
XFILL_8_NAND2X1_81 gnd vdd FILL
XFILL_30_DFFSR_154 gnd vdd FILL
XFILL_3_INVX8_4 gnd vdd FILL
XFILL_8_NAND2X1_92 gnd vdd FILL
XFILL_30_DFFSR_165 gnd vdd FILL
XFILL_16_INVX8_2 gnd vdd FILL
XFILL_30_DFFSR_176 gnd vdd FILL
XFILL_30_DFFSR_187 gnd vdd FILL
XFILL_16_CLKBUF1_12 gnd vdd FILL
XFILL_30_DFFSR_198 gnd vdd FILL
XFILL_34_DFFSR_120 gnd vdd FILL
XFILL_16_CLKBUF1_23 gnd vdd FILL
XFILL_34_DFFSR_131 gnd vdd FILL
XFILL_16_CLKBUF1_34 gnd vdd FILL
XFILL_34_DFFSR_142 gnd vdd FILL
XFILL_11_AOI21X1_20 gnd vdd FILL
XFILL_34_DFFSR_153 gnd vdd FILL
XFILL_11_AOI21X1_31 gnd vdd FILL
XFILL_34_DFFSR_164 gnd vdd FILL
XFILL_34_DFFSR_175 gnd vdd FILL
XFILL_11_AOI21X1_42 gnd vdd FILL
XFILL_34_DFFSR_186 gnd vdd FILL
XFILL_11_AOI21X1_53 gnd vdd FILL
XFILL_20_DFFSR_4 gnd vdd FILL
XFILL_34_DFFSR_197 gnd vdd FILL
XFILL_11_AOI21X1_64 gnd vdd FILL
XFILL_11_AOI21X1_75 gnd vdd FILL
XFILL_38_DFFSR_130 gnd vdd FILL
XFILL_38_DFFSR_141 gnd vdd FILL
XFILL_38_DFFSR_152 gnd vdd FILL
XFILL_58_DFFSR_2 gnd vdd FILL
XFILL_38_DFFSR_163 gnd vdd FILL
XFILL_38_DFFSR_174 gnd vdd FILL
XFILL_2_INVX1_18 gnd vdd FILL
XFILL_30_NOR3X1_10 gnd vdd FILL
XFILL_2_INVX1_29 gnd vdd FILL
XFILL_38_DFFSR_185 gnd vdd FILL
XFILL_30_NOR3X1_21 gnd vdd FILL
XFILL_38_DFFSR_196 gnd vdd FILL
XFILL_30_NOR3X1_32 gnd vdd FILL
XFILL_30_NOR3X1_43 gnd vdd FILL
XFILL_80_DFFSR_210 gnd vdd FILL
XFILL_80_DFFSR_221 gnd vdd FILL
XFILL_80_DFFSR_232 gnd vdd FILL
XFILL_80_DFFSR_243 gnd vdd FILL
XFILL_80_DFFSR_254 gnd vdd FILL
XFILL_80_DFFSR_265 gnd vdd FILL
XFILL_16_DFFSR_109 gnd vdd FILL
XFILL_84_DFFSR_220 gnd vdd FILL
XFILL_0_BUFX4_16 gnd vdd FILL
XFILL_11_AOI21X1_5 gnd vdd FILL
XFILL_84_DFFSR_231 gnd vdd FILL
XFILL_0_BUFX4_27 gnd vdd FILL
XFILL_84_DFFSR_242 gnd vdd FILL
XFILL_42_DFFSR_8 gnd vdd FILL
XFILL_37_6_1 gnd vdd FILL
XFILL_84_DFFSR_253 gnd vdd FILL
XFILL_36_1_0 gnd vdd FILL
XFILL_0_BUFX4_38 gnd vdd FILL
XFILL_84_DFFSR_264 gnd vdd FILL
XFILL_0_BUFX4_49 gnd vdd FILL
XFILL_84_DFFSR_275 gnd vdd FILL
XFILL_6_CLKBUF1_40 gnd vdd FILL
XFILL_14_MUX2X1_103 gnd vdd FILL
XFILL_14_MUX2X1_114 gnd vdd FILL
XFILL_14_MUX2X1_125 gnd vdd FILL
XFILL_14_MUX2X1_136 gnd vdd FILL
XFILL_15_AOI21X1_4 gnd vdd FILL
XFILL_0_INVX1_170 gnd vdd FILL
XFILL_0_INVX1_181 gnd vdd FILL
XFILL_14_MUX2X1_147 gnd vdd FILL
XFILL_14_MUX2X1_158 gnd vdd FILL
XFILL_57_DFFSR_19 gnd vdd FILL
XFILL_1_AOI21X1_70 gnd vdd FILL
XFILL_14_MUX2X1_169 gnd vdd FILL
XFILL_0_INVX1_192 gnd vdd FILL
XFILL_1_AOI21X1_81 gnd vdd FILL
XFILL_28_10 gnd vdd FILL
XFILL_11_OAI22X1_50 gnd vdd FILL
XFILL_15_OAI21X1_30 gnd vdd FILL
XFILL_15_OAI21X1_41 gnd vdd FILL
XFILL_20_5_1 gnd vdd FILL
XFILL_4_INVX1_180 gnd vdd FILL
XFILL_4_INVX1_191 gnd vdd FILL
XFILL_4_NOR2X1_180 gnd vdd FILL
XFILL_4_NOR2X1_191 gnd vdd FILL
XFILL_66_DFFSR_209 gnd vdd FILL
XFILL_26_DFFSR_18 gnd vdd FILL
XFILL_26_DFFSR_29 gnd vdd FILL
XFILL_66_DFFSR_17 gnd vdd FILL
XFILL_66_DFFSR_28 gnd vdd FILL
XFILL_66_DFFSR_39 gnd vdd FILL
XFILL_21_MUX2X1_160 gnd vdd FILL
XFILL_21_MUX2X1_171 gnd vdd FILL
XNAND3X1_16 NAND3X1_16/A NAND3X1_16/B NAND3X1_16/C gnd INVX1_129/A vdd NAND3X1
XFILL_21_MUX2X1_182 gnd vdd FILL
XFILL_4_MUX2X1_120 gnd vdd FILL
XFILL_21_MUX2X1_193 gnd vdd FILL
XNAND3X1_27 BUFX2_8/A OAI21X1_33/Y OAI21X1_35/Y gnd AOI22X1_1/A vdd NAND3X1
XFILL_4_MUX2X1_131 gnd vdd FILL
XFILL_4_MUX2X1_142 gnd vdd FILL
XNAND3X1_38 INVX1_134/Y INVX1_137/A INVX1_57/A gnd NAND3X1_38/Y vdd NAND3X1
XFILL_4_MUX2X1_153 gnd vdd FILL
XNAND3X1_49 NOR3X1_9/A DFFSR_199/D AND2X2_6/B gnd NOR3X1_6/B vdd NAND3X1
XFILL_9_DFFSR_19 gnd vdd FILL
XFILL_4_BUFX4_7 gnd vdd FILL
XFILL_4_MUX2X1_164 gnd vdd FILL
XFILL_4_MUX2X1_175 gnd vdd FILL
XFILL_7_NAND3X1_108 gnd vdd FILL
XFILL_4_MUX2X1_186 gnd vdd FILL
XFILL_35_DFFSR_16 gnd vdd FILL
XFILL_7_NAND3X1_119 gnd vdd FILL
XFILL_35_DFFSR_27 gnd vdd FILL
XFILL_35_DFFSR_38 gnd vdd FILL
XNOR2X1_16 NOR2X1_16/A NOR2X1_16/B gnd NOR2X1_16/Y vdd NOR2X1
XNOR2X1_27 NOR2X1_27/A OR2X2_1/A gnd NOR2X1_28/B vdd NOR2X1
XFILL_35_DFFSR_49 gnd vdd FILL
XFILL_28_6_1 gnd vdd FILL
XFILL_3_6_1 gnd vdd FILL
XNOR2X1_38 NOR3X1_9/C NOR2X1_44/B gnd NOR2X1_38/Y vdd NOR2X1
XNOR2X1_49 NOR2X1_49/A NOR2X1_49/B gnd NOR2X1_49/Y vdd NOR2X1
XFILL_2_1_0 gnd vdd FILL
XFILL_51_DFFSR_220 gnd vdd FILL
XFILL_27_1_0 gnd vdd FILL
XFILL_51_DFFSR_231 gnd vdd FILL
XFILL_51_DFFSR_242 gnd vdd FILL
XFILL_51_DFFSR_253 gnd vdd FILL
XFILL_75_DFFSR_15 gnd vdd FILL
XFILL_75_DFFSR_26 gnd vdd FILL
XFILL_51_DFFSR_264 gnd vdd FILL
XFILL_51_DFFSR_275 gnd vdd FILL
XFILL_75_DFFSR_37 gnd vdd FILL
XFILL_75_DFFSR_48 gnd vdd FILL
XFILL_18_MUX2X1_5 gnd vdd FILL
XFILL_75_DFFSR_59 gnd vdd FILL
XFILL_55_DFFSR_230 gnd vdd FILL
XFILL_55_DFFSR_241 gnd vdd FILL
XFILL_55_DFFSR_252 gnd vdd FILL
XFILL_11_NAND3X1_110 gnd vdd FILL
XFILL_11_NAND3X1_121 gnd vdd FILL
XFILL_10_CLKBUF1_4 gnd vdd FILL
XFILL_11_NAND3X1_132 gnd vdd FILL
XFILL_55_DFFSR_263 gnd vdd FILL
XFILL_55_DFFSR_274 gnd vdd FILL
XFILL_10_NAND2X1_19 gnd vdd FILL
XFILL_11_5_1 gnd vdd FILL
XFILL_9_BUFX4_60 gnd vdd FILL
XFILL_44_DFFSR_14 gnd vdd FILL
XFILL_0_BUFX2_3 gnd vdd FILL
XFILL_9_BUFX4_71 gnd vdd FILL
XFILL_44_DFFSR_25 gnd vdd FILL
XFILL_82_DFFSR_130 gnd vdd FILL
XFILL_10_0_0 gnd vdd FILL
XFILL_9_BUFX4_82 gnd vdd FILL
XFILL_9_BUFX4_93 gnd vdd FILL
XFILL_44_DFFSR_36 gnd vdd FILL
XFILL_59_DFFSR_240 gnd vdd FILL
XFILL_82_DFFSR_141 gnd vdd FILL
XFILL_44_DFFSR_47 gnd vdd FILL
XFILL_82_DFFSR_152 gnd vdd FILL
XFILL_44_DFFSR_58 gnd vdd FILL
XFILL_59_DFFSR_251 gnd vdd FILL
XFILL_59_DFFSR_262 gnd vdd FILL
XFILL_44_DFFSR_69 gnd vdd FILL
XFILL_82_DFFSR_163 gnd vdd FILL
XFILL_82_DFFSR_174 gnd vdd FILL
XFILL_14_CLKBUF1_3 gnd vdd FILL
XFILL_2_DFFSR_200 gnd vdd FILL
XFILL_59_DFFSR_273 gnd vdd FILL
XFILL_82_DFFSR_185 gnd vdd FILL
XFILL_84_DFFSR_13 gnd vdd FILL
XFILL_2_DFFSR_211 gnd vdd FILL
XFILL_82_DFFSR_196 gnd vdd FILL
XFILL_2_DFFSR_222 gnd vdd FILL
XFILL_84_DFFSR_24 gnd vdd FILL
XFILL_7_NAND3X1_12 gnd vdd FILL
XFILL_33_DFFSR_209 gnd vdd FILL
XFILL_84_DFFSR_35 gnd vdd FILL
XFILL_2_DFFSR_233 gnd vdd FILL
XFILL_7_NAND3X1_23 gnd vdd FILL
XFILL_86_DFFSR_140 gnd vdd FILL
XFILL_2_DFFSR_244 gnd vdd FILL
XFILL_84_DFFSR_46 gnd vdd FILL
XFILL_7_NAND3X1_34 gnd vdd FILL
XFILL_2_NAND3X1_104 gnd vdd FILL
XFILL_13_DFFSR_13 gnd vdd FILL
XFILL_84_DFFSR_57 gnd vdd FILL
XFILL_86_DFFSR_151 gnd vdd FILL
XFILL_2_DFFSR_255 gnd vdd FILL
XFILL_2_NAND3X1_115 gnd vdd FILL
XFILL_7_NAND3X1_45 gnd vdd FILL
XFILL_86_DFFSR_162 gnd vdd FILL
XFILL_84_DFFSR_68 gnd vdd FILL
XFILL_13_DFFSR_24 gnd vdd FILL
XFILL_7_NAND3X1_56 gnd vdd FILL
XFILL_2_NAND3X1_126 gnd vdd FILL
XFILL_2_DFFSR_266 gnd vdd FILL
XFILL_13_DFFSR_35 gnd vdd FILL
XFILL_86_DFFSR_173 gnd vdd FILL
XFILL_84_DFFSR_79 gnd vdd FILL
XFILL_7_NAND3X1_67 gnd vdd FILL
XFILL_18_CLKBUF1_2 gnd vdd FILL
XFILL_86_DFFSR_184 gnd vdd FILL
XFILL_7_NAND3X1_78 gnd vdd FILL
XFILL_6_DFFSR_210 gnd vdd FILL
XFILL_13_DFFSR_46 gnd vdd FILL
XFILL_86_DFFSR_195 gnd vdd FILL
XFILL_60_DFFSR_109 gnd vdd FILL
XFILL_13_DFFSR_57 gnd vdd FILL
XFILL_7_NAND3X1_89 gnd vdd FILL
XFILL_37_DFFSR_208 gnd vdd FILL
XFILL_13_DFFSR_68 gnd vdd FILL
XFILL_6_DFFSR_221 gnd vdd FILL
XFILL_37_DFFSR_219 gnd vdd FILL
XFILL_13_DFFSR_79 gnd vdd FILL
XFILL_6_DFFSR_232 gnd vdd FILL
XFILL_6_DFFSR_243 gnd vdd FILL
XFILL_6_DFFSR_254 gnd vdd FILL
XFILL_53_DFFSR_12 gnd vdd FILL
XFILL_53_DFFSR_23 gnd vdd FILL
XFILL_6_DFFSR_265 gnd vdd FILL
XFILL_53_DFFSR_34 gnd vdd FILL
XFILL_24_NOR3X1_9 gnd vdd FILL
XFILL_53_DFFSR_45 gnd vdd FILL
XFILL_53_DFFSR_56 gnd vdd FILL
XFILL_64_DFFSR_108 gnd vdd FILL
XFILL_53_DFFSR_67 gnd vdd FILL
XFILL_64_DFFSR_119 gnd vdd FILL
XFILL_53_DFFSR_78 gnd vdd FILL
XFILL_53_DFFSR_89 gnd vdd FILL
XFILL_14_AOI21X1_19 gnd vdd FILL
XFILL_19_6_1 gnd vdd FILL
XFILL_0_NAND2X1_14 gnd vdd FILL
XMUX2X1_12 MUX2X1_9/A INVX1_26/Y MUX2X1_14/S gnd DFFSR_33/D vdd MUX2X1
XMUX2X1_23 BUFX4_63/Y INVX1_37/Y NOR2X1_9/B gnd MUX2X1_23/Y vdd MUX2X1
XFILL_0_NAND2X1_25 gnd vdd FILL
XMUX2X1_34 BUFX4_77/Y INVX1_48/Y NOR2X1_20/Y gnd MUX2X1_34/Y vdd MUX2X1
XFILL_18_1_0 gnd vdd FILL
XFILL_0_NAND2X1_36 gnd vdd FILL
XFILL_24_DFFSR_5 gnd vdd FILL
XNOR2X1_106 OAI21X1_30/Y OAI22X1_46/Y gnd NOR2X1_106/Y vdd NOR2X1
XMUX2X1_45 INVX1_59/Y MUX2X1_4/B NAND2X1_7/Y gnd MUX2X1_45/Y vdd MUX2X1
XFILL_0_NAND2X1_47 gnd vdd FILL
XFILL_68_DFFSR_107 gnd vdd FILL
XFILL_22_DFFSR_11 gnd vdd FILL
XMUX2X1_56 INVX1_70/Y BUFX4_71/Y NAND2X1_9/Y gnd MUX2X1_56/Y vdd MUX2X1
XNOR2X1_117 OAI21X1_47/A NOR3X1_48/Y gnd DFFSR_199/D vdd NOR2X1
XFILL_81_DFFSR_6 gnd vdd FILL
XNOR2X1_128 NOR2X1_25/A INVX4_1/Y gnd NOR2X1_128/Y vdd NOR2X1
XFILL_0_NAND2X1_58 gnd vdd FILL
XFILL_22_DFFSR_22 gnd vdd FILL
XFILL_68_DFFSR_118 gnd vdd FILL
XFILL_0_NAND2X1_69 gnd vdd FILL
XFILL_68_DFFSR_129 gnd vdd FILL
XFILL_22_DFFSR_33 gnd vdd FILL
XMUX2X1_67 INVX1_81/Y BUFX4_86/Y MUX2X1_71/S gnd MUX2X1_67/Y vdd MUX2X1
XMUX2X1_78 BUFX4_96/Y INVX1_92/Y NOR2X1_26/B gnd MUX2X1_78/Y vdd MUX2X1
XNOR2X1_139 NOR2X1_20/A INVX4_1/Y gnd NOR2X1_139/Y vdd NOR2X1
XFILL_22_DFFSR_44 gnd vdd FILL
XFILL_22_DFFSR_55 gnd vdd FILL
XMUX2X1_89 MUX2X1_89/A BUFX4_75/Y MUX2X1_91/S gnd MUX2X1_89/Y vdd MUX2X1
XFILL_61_4_1 gnd vdd FILL
XFILL_11_OAI21X1_8 gnd vdd FILL
XFILL_0_INVX2_3 gnd vdd FILL
XFILL_22_DFFSR_66 gnd vdd FILL
XFILL_22_DFFSR_77 gnd vdd FILL
XFILL_22_DFFSR_88 gnd vdd FILL
XFILL_22_DFFSR_99 gnd vdd FILL
XFILL_62_DFFSR_10 gnd vdd FILL
XFILL_23_5 gnd vdd FILL
XFILL_62_DFFSR_21 gnd vdd FILL
XFILL_62_DFFSR_32 gnd vdd FILL
XFILL_62_DFFSR_43 gnd vdd FILL
XFILL_16_4 gnd vdd FILL
XFILL_22_DFFSR_230 gnd vdd FILL
XFILL_62_DFFSR_54 gnd vdd FILL
XFILL_3_AOI22X1_4 gnd vdd FILL
XFILL_15_OAI21X1_7 gnd vdd FILL
XFILL_22_DFFSR_241 gnd vdd FILL
XFILL_62_DFFSR_65 gnd vdd FILL
XFILL_22_DFFSR_252 gnd vdd FILL
XFILL_62_DFFSR_76 gnd vdd FILL
XFILL_62_DFFSR_87 gnd vdd FILL
XFILL_22_DFFSR_263 gnd vdd FILL
XFILL_22_DFFSR_274 gnd vdd FILL
XFILL_62_DFFSR_98 gnd vdd FILL
XFILL_3_INVX1_203 gnd vdd FILL
XFILL_3_INVX1_214 gnd vdd FILL
XFILL_26_CLKBUF1_13 gnd vdd FILL
XDFFSR_4 DFFSR_4/Q DFFSR_4/CLK DFFSR_4/R vdd DFFSR_4/D gnd vdd DFFSR
XFILL_5_DFFSR_12 gnd vdd FILL
XFILL_26_CLKBUF1_24 gnd vdd FILL
XFILL_3_INVX1_225 gnd vdd FILL
XFILL_26_CLKBUF1_35 gnd vdd FILL
XFILL_7_AOI22X1_3 gnd vdd FILL
XFILL_5_DFFSR_23 gnd vdd FILL
XFILL_5_DFFSR_34 gnd vdd FILL
XFILL_31_DFFSR_20 gnd vdd FILL
XFILL_5_DFFSR_45 gnd vdd FILL
XFILL_26_DFFSR_240 gnd vdd FILL
XFILL_46_DFFSR_9 gnd vdd FILL
XFILL_5_DFFSR_56 gnd vdd FILL
XFILL_26_DFFSR_251 gnd vdd FILL
XFILL_26_DFFSR_262 gnd vdd FILL
XFILL_31_DFFSR_31 gnd vdd FILL
XFILL_5_DFFSR_67 gnd vdd FILL
XFILL_31_DFFSR_42 gnd vdd FILL
XFILL_5_DFFSR_78 gnd vdd FILL
XFILL_7_INVX1_202 gnd vdd FILL
XFILL_31_DFFSR_53 gnd vdd FILL
XFILL_26_DFFSR_273 gnd vdd FILL
XFILL_9_CLKBUF1_17 gnd vdd FILL
XFILL_9_CLKBUF1_28 gnd vdd FILL
XFILL_5_DFFSR_89 gnd vdd FILL
XFILL_23_MUX2X1_18 gnd vdd FILL
XFILL_31_DFFSR_64 gnd vdd FILL
XFILL_23_MUX2X1_29 gnd vdd FILL
XFILL_7_INVX1_213 gnd vdd FILL
XFILL_31_DFFSR_75 gnd vdd FILL
XFILL_9_CLKBUF1_39 gnd vdd FILL
XFILL_7_INVX1_224 gnd vdd FILL
XFILL_31_DFFSR_86 gnd vdd FILL
XFILL_4_AOI21X1_14 gnd vdd FILL
XFILL_53_DFFSR_140 gnd vdd FILL
XFILL_4_AOI21X1_25 gnd vdd FILL
XFILL_31_DFFSR_97 gnd vdd FILL
XFILL_4_AOI21X1_36 gnd vdd FILL
XFILL_53_DFFSR_151 gnd vdd FILL
XFILL_4_AOI21X1_47 gnd vdd FILL
XFILL_71_DFFSR_30 gnd vdd FILL
XFILL_53_DFFSR_162 gnd vdd FILL
XFILL_4_AOI21X1_58 gnd vdd FILL
XFILL_53_DFFSR_173 gnd vdd FILL
XFILL_71_DFFSR_41 gnd vdd FILL
XFILL_14_OAI22X1_16 gnd vdd FILL
XFILL_53_DFFSR_184 gnd vdd FILL
XFILL_4_AOI21X1_69 gnd vdd FILL
XFILL_14_OAI22X1_27 gnd vdd FILL
XFILL_71_DFFSR_52 gnd vdd FILL
XFILL_71_DFFSR_63 gnd vdd FILL
XFILL_14_OAI22X1_38 gnd vdd FILL
XINVX1_19 INVX1_19/A gnd MUX2X1_6/A vdd INVX1
XFILL_53_DFFSR_195 gnd vdd FILL
XFILL_71_DFFSR_74 gnd vdd FILL
XFILL_7_NOR2X1_102 gnd vdd FILL
XFILL_71_DFFSR_85 gnd vdd FILL
XFILL_14_OAI22X1_49 gnd vdd FILL
XFILL_7_NOR2X1_113 gnd vdd FILL
XFILL_7_NOR2X1_124 gnd vdd FILL
XFILL_71_DFFSR_96 gnd vdd FILL
XFILL_57_DFFSR_150 gnd vdd FILL
XFILL_7_NOR2X1_135 gnd vdd FILL
XFILL_7_NOR2X1_146 gnd vdd FILL
XFILL_57_DFFSR_161 gnd vdd FILL
XFILL_7_NOR2X1_157 gnd vdd FILL
XFILL_57_DFFSR_172 gnd vdd FILL
XFILL_57_DFFSR_183 gnd vdd FILL
XFILL_7_NOR2X1_168 gnd vdd FILL
XFILL_7_NOR2X1_179 gnd vdd FILL
XFILL_57_DFFSR_194 gnd vdd FILL
XFILL_0_DFFSR_110 gnd vdd FILL
XFILL_31_DFFSR_108 gnd vdd FILL
XNAND2X1_60 NOR2X1_59/Y NOR2X1_58/Y gnd NOR3X1_11/B vdd NAND2X1
XFILL_0_DFFSR_121 gnd vdd FILL
XFILL_40_DFFSR_40 gnd vdd FILL
XFILL_0_DFFSR_132 gnd vdd FILL
XFILL_13_NAND3X1_70 gnd vdd FILL
XFILL_31_DFFSR_119 gnd vdd FILL
XNAND2X1_71 BUFX4_103/Y AND2X2_3/Y gnd OAI22X1_36/D vdd NAND2X1
XFILL_11_NOR3X1_4 gnd vdd FILL
XFILL_13_NAND3X1_81 gnd vdd FILL
XNAND2X1_82 INVX2_4/A INVX2_5/A gnd NOR2X1_24/A vdd NAND2X1
XFILL_40_DFFSR_51 gnd vdd FILL
XFILL_0_DFFSR_143 gnd vdd FILL
XFILL_13_NAND3X1_92 gnd vdd FILL
XNAND2X1_93 NAND3X1_33/Y OAI21X1_41/Y gnd DFFSR_1/D vdd NAND2X1
XFILL_0_DFFSR_154 gnd vdd FILL
XFILL_40_DFFSR_62 gnd vdd FILL
XFILL_0_DFFSR_165 gnd vdd FILL
XFILL_40_DFFSR_73 gnd vdd FILL
XFILL_40_DFFSR_84 gnd vdd FILL
XFILL_0_DFFSR_176 gnd vdd FILL
XFILL_40_DFFSR_95 gnd vdd FILL
XFILL_0_DFFSR_187 gnd vdd FILL
XFILL_0_DFFSR_198 gnd vdd FILL
XFILL_35_DFFSR_107 gnd vdd FILL
XFILL_4_DFFSR_120 gnd vdd FILL
XFILL_4_DFFSR_131 gnd vdd FILL
XFILL_52_4_1 gnd vdd FILL
XFILL_35_DFFSR_118 gnd vdd FILL
XFILL_4_DFFSR_142 gnd vdd FILL
XFILL_35_DFFSR_129 gnd vdd FILL
XFILL_80_DFFSR_50 gnd vdd FILL
XFILL_4_DFFSR_153 gnd vdd FILL
XFILL_80_DFFSR_61 gnd vdd FILL
XFILL_80_DFFSR_72 gnd vdd FILL
XFILL_4_DFFSR_164 gnd vdd FILL
XFILL_80_DFFSR_83 gnd vdd FILL
XFILL_4_DFFSR_175 gnd vdd FILL
XFILL_4_DFFSR_186 gnd vdd FILL
XFILL_80_DFFSR_94 gnd vdd FILL
XFILL_4_DFFSR_197 gnd vdd FILL
XFILL_7_MUX2X1_108 gnd vdd FILL
XFILL_39_DFFSR_106 gnd vdd FILL
XFILL_7_MUX2X1_119 gnd vdd FILL
XFILL_8_DFFSR_130 gnd vdd FILL
XFILL_39_DFFSR_117 gnd vdd FILL
XFILL_39_DFFSR_128 gnd vdd FILL
XFILL_8_DFFSR_141 gnd vdd FILL
XFILL_39_DFFSR_139 gnd vdd FILL
XFILL_8_DFFSR_152 gnd vdd FILL
XFILL_4_OAI22X1_11 gnd vdd FILL
XFILL_8_BUFX4_8 gnd vdd FILL
XFILL_12_MUX2X1_50 gnd vdd FILL
XFILL_8_DFFSR_163 gnd vdd FILL
XFILL_12_MUX2X1_61 gnd vdd FILL
XFILL_8_DFFSR_174 gnd vdd FILL
XFILL_0_NOR3X1_10 gnd vdd FILL
XFILL_20_NOR3X1_2 gnd vdd FILL
XFILL_4_OAI22X1_22 gnd vdd FILL
XFILL_12_MUX2X1_72 gnd vdd FILL
XFILL_12_MUX2X1_83 gnd vdd FILL
XFILL_4_OAI22X1_33 gnd vdd FILL
XFILL_8_DFFSR_185 gnd vdd FILL
XFILL_12_MUX2X1_94 gnd vdd FILL
XFILL_4_OAI22X1_44 gnd vdd FILL
XFILL_0_NOR3X1_21 gnd vdd FILL
XFILL_8_DFFSR_196 gnd vdd FILL
XFILL_0_NOR3X1_32 gnd vdd FILL
XFILL_31_NOR3X1_19 gnd vdd FILL
XFILL_8_OAI21X1_13 gnd vdd FILL
XFILL_0_NOR3X1_43 gnd vdd FILL
XFILL_8_OAI21X1_24 gnd vdd FILL
XFILL_8_OAI21X1_35 gnd vdd FILL
XFILL_81_DFFSR_208 gnd vdd FILL
XFILL_81_DFFSR_219 gnd vdd FILL
XFILL_8_OAI21X1_46 gnd vdd FILL
XFILL_16_MUX2X1_60 gnd vdd FILL
XFILL_16_MUX2X1_71 gnd vdd FILL
XFILL_16_MUX2X1_82 gnd vdd FILL
XFILL_4_NOR3X1_20 gnd vdd FILL
XFILL_16_MUX2X1_93 gnd vdd FILL
XFILL_4_NOR3X1_31 gnd vdd FILL
XFILL_4_NOR3X1_42 gnd vdd FILL
XFILL_85_DFFSR_207 gnd vdd FILL
XFILL_1_NOR2X1_202 gnd vdd FILL
XFILL_85_DFFSR_218 gnd vdd FILL
XFILL_20_DFFSR_140 gnd vdd FILL
XFILL_85_DFFSR_229 gnd vdd FILL
XFILL_20_DFFSR_151 gnd vdd FILL
XFILL_20_DFFSR_162 gnd vdd FILL
XFILL_3_NOR3X1_3 gnd vdd FILL
XFILL_20_DFFSR_173 gnd vdd FILL
XFILL_8_NOR3X1_30 gnd vdd FILL
XFILL_20_DFFSR_184 gnd vdd FILL
XFILL_1_INVX1_102 gnd vdd FILL
XFILL_59_0_0 gnd vdd FILL
XFILL_1_INVX1_113 gnd vdd FILL
XFILL_8_NOR3X1_41 gnd vdd FILL
XFILL_8_NOR3X1_52 gnd vdd FILL
XFILL_1_INVX1_124 gnd vdd FILL
XFILL_20_DFFSR_195 gnd vdd FILL
XFILL_15_CLKBUF1_20 gnd vdd FILL
XFILL_1_INVX1_135 gnd vdd FILL
XFILL_4_BUFX2_4 gnd vdd FILL
XFILL_15_CLKBUF1_31 gnd vdd FILL
XFILL_1_INVX1_146 gnd vdd FILL
XFILL_15_CLKBUF1_42 gnd vdd FILL
XFILL_1_INVX1_157 gnd vdd FILL
XFILL_1_INVX1_168 gnd vdd FILL
XFILL_24_DFFSR_150 gnd vdd FILL
XFILL_24_DFFSR_161 gnd vdd FILL
XFILL_1_INVX1_179 gnd vdd FILL
XFILL_24_DFFSR_172 gnd vdd FILL
XFILL_8_NAND3X1_109 gnd vdd FILL
XFILL_24_DFFSR_183 gnd vdd FILL
XFILL_5_INVX1_101 gnd vdd FILL
XFILL_10_AOI21X1_50 gnd vdd FILL
XFILL_5_INVX1_112 gnd vdd FILL
XFILL_24_DFFSR_194 gnd vdd FILL
XFILL_5_INVX1_123 gnd vdd FILL
XFILL_10_AOI21X1_61 gnd vdd FILL
XFILL_10_AOI21X1_72 gnd vdd FILL
XFILL_5_INVX1_134 gnd vdd FILL
XFILL_5_INVX1_145 gnd vdd FILL
XFILL_63_DFFSR_3 gnd vdd FILL
XFILL_5_INVX1_156 gnd vdd FILL
XFILL_1_DFFSR_60 gnd vdd FILL
XFILL_5_INVX1_167 gnd vdd FILL
XFILL_1_DFFSR_71 gnd vdd FILL
XFILL_28_DFFSR_160 gnd vdd FILL
XFILL_43_4_1 gnd vdd FILL
XFILL_5_INVX1_178 gnd vdd FILL
XFILL_1_DFFSR_82 gnd vdd FILL
XFILL_5_INVX1_189 gnd vdd FILL
XFILL_28_DFFSR_171 gnd vdd FILL
XFILL_1_DFFSR_93 gnd vdd FILL
XFILL_28_DFFSR_182 gnd vdd FILL
XFILL_28_DFFSR_193 gnd vdd FILL
XFILL_20_NOR3X1_40 gnd vdd FILL
XFILL_20_NOR3X1_51 gnd vdd FILL
XFILL_12_NAND3X1_100 gnd vdd FILL
XFILL_70_DFFSR_240 gnd vdd FILL
XFILL_70_DFFSR_251 gnd vdd FILL
XFILL_12_NAND3X1_111 gnd vdd FILL
XFILL_12_NAND3X1_122 gnd vdd FILL
XFILL_70_DFFSR_262 gnd vdd FILL
XFILL_70_DFFSR_273 gnd vdd FILL
XFILL_24_NOR3X1_50 gnd vdd FILL
XFILL_3_OAI22X1_7 gnd vdd FILL
XFILL_74_DFFSR_250 gnd vdd FILL
XFILL_74_DFFSR_261 gnd vdd FILL
XFILL_28_DFFSR_6 gnd vdd FILL
XFILL_74_DFFSR_272 gnd vdd FILL
XFILL_85_DFFSR_7 gnd vdd FILL
XFILL_13_MUX2X1_100 gnd vdd FILL
XFILL_13_MUX2X1_111 gnd vdd FILL
XFILL_13_MUX2X1_122 gnd vdd FILL
XFILL_7_OAI22X1_6 gnd vdd FILL
XFILL_4_INVX2_4 gnd vdd FILL
XFILL_13_MUX2X1_133 gnd vdd FILL
XFILL_13_MUX2X1_144 gnd vdd FILL
XFILL_3_NAND3X1_105 gnd vdd FILL
XFILL_3_NAND3X1_116 gnd vdd FILL
XFILL_13_MUX2X1_155 gnd vdd FILL
XFILL_78_DFFSR_260 gnd vdd FILL
XFILL_3_NAND3X1_127 gnd vdd FILL
XFILL_78_DFFSR_271 gnd vdd FILL
XFILL_33_CLKBUF1_1 gnd vdd FILL
XFILL_13_MUX2X1_166 gnd vdd FILL
XFILL_13_MUX2X1_177 gnd vdd FILL
XFILL_13_MUX2X1_188 gnd vdd FILL
XFILL_52_DFFSR_207 gnd vdd FILL
XFILL_52_DFFSR_218 gnd vdd FILL
XFILL_52_DFFSR_229 gnd vdd FILL
XFILL_2_INVX1_2 gnd vdd FILL
XFILL_56_DFFSR_206 gnd vdd FILL
XFILL_56_DFFSR_217 gnd vdd FILL
XFILL_56_DFFSR_228 gnd vdd FILL
XFILL_56_DFFSR_239 gnd vdd FILL
XFILL_83_DFFSR_106 gnd vdd FILL
XFILL_34_4_1 gnd vdd FILL
XFILL_83_DFFSR_117 gnd vdd FILL
XFILL_83_DFFSR_128 gnd vdd FILL
XFILL_83_DFFSR_139 gnd vdd FILL
XFILL_21_2 gnd vdd FILL
XFILL_87_DFFSR_105 gnd vdd FILL
XFILL_20_MUX2X1_190 gnd vdd FILL
XFILL_14_1 gnd vdd FILL
XFILL_0_NAND3X1_9 gnd vdd FILL
XFILL_3_DFFSR_209 gnd vdd FILL
XFILL_87_DFFSR_116 gnd vdd FILL
XFILL_14_BUFX4_10 gnd vdd FILL
XFILL_87_DFFSR_127 gnd vdd FILL
XFILL_87_DFFSR_138 gnd vdd FILL
XFILL_3_MUX2X1_150 gnd vdd FILL
XFILL_14_BUFX4_21 gnd vdd FILL
XFILL_3_MUX2X1_161 gnd vdd FILL
XFILL_87_DFFSR_149 gnd vdd FILL
XFILL_14_BUFX4_32 gnd vdd FILL
XFILL_14_BUFX4_43 gnd vdd FILL
XFILL_3_MUX2X1_172 gnd vdd FILL
XDFFSR_200 INVX1_99/A DFFSR_57/CLK BUFX4_21/Y vdd MUX2X1_86/Y gnd vdd DFFSR
XFILL_14_BUFX4_54 gnd vdd FILL
XFILL_3_MUX2X1_183 gnd vdd FILL
XDFFSR_211 INVX1_86/A DFFSR_45/CLK DFFSR_57/R vdd MUX2X1_73/Y gnd vdd DFFSR
XFILL_14_BUFX4_65 gnd vdd FILL
XFILL_3_MUX2X1_194 gnd vdd FILL
XFILL_7_DFFSR_208 gnd vdd FILL
XFILL_14_BUFX4_76 gnd vdd FILL
XDFFSR_222 INVX1_80/A DFFSR_4/CLK DFFSR_4/R vdd MUX2X1_66/Y gnd vdd DFFSR
XFILL_4_NAND3X1_8 gnd vdd FILL
XFILL_7_DFFSR_219 gnd vdd FILL
XDFFSR_233 INVX1_64/A DFFSR_58/CLK DFFSR_23/R vdd MUX2X1_51/Y gnd vdd DFFSR
XFILL_14_BUFX4_87 gnd vdd FILL
XDFFSR_244 INVX1_58/A CLKBUF1_34/Y BUFX4_23/Y vdd MUX2X1_44/Y gnd vdd DFFSR
XFILL_14_BUFX4_98 gnd vdd FILL
XDFFSR_255 INVX1_43/A DFFSR_5/CLK DFFSR_5/R vdd MUX2X1_30/Y gnd vdd DFFSR
XDFFSR_266 NOR2X1_12/A DFFSR_9/CLK BUFX4_54/Y vdd DFFSR_266/D gnd vdd DFFSR
XFILL_41_DFFSR_250 gnd vdd FILL
XFILL_41_DFFSR_261 gnd vdd FILL
XFILL_41_DFFSR_272 gnd vdd FILL
XFILL_8_NAND3X1_7 gnd vdd FILL
XFILL_45_DFFSR_260 gnd vdd FILL
XFILL_45_DFFSR_271 gnd vdd FILL
XFILL_9_AND2X2_3 gnd vdd FILL
XFILL_72_DFFSR_160 gnd vdd FILL
XFILL_49_DFFSR_270 gnd vdd FILL
XFILL_72_DFFSR_171 gnd vdd FILL
XFILL_72_DFFSR_182 gnd vdd FILL
XFILL_72_DFFSR_19 gnd vdd FILL
XFILL_72_DFFSR_193 gnd vdd FILL
XFILL_23_DFFSR_206 gnd vdd FILL
XFILL_6_NAND3X1_20 gnd vdd FILL
XFILL_23_DFFSR_217 gnd vdd FILL
XFILL_23_DFFSR_228 gnd vdd FILL
XFILL_6_NAND3X1_31 gnd vdd FILL
XFILL_23_DFFSR_239 gnd vdd FILL
XFILL_15_MUX2X1_9 gnd vdd FILL
XFILL_6_NAND3X1_42 gnd vdd FILL
XFILL_6_NAND3X1_53 gnd vdd FILL
XFILL_0_4_1 gnd vdd FILL
XFILL_25_4_1 gnd vdd FILL
XFILL_76_DFFSR_170 gnd vdd FILL
XFILL_6_NAND3X1_64 gnd vdd FILL
XFILL_6_NAND3X1_75 gnd vdd FILL
XFILL_76_DFFSR_181 gnd vdd FILL
XFILL_6_BUFX4_20 gnd vdd FILL
XFILL_6_NAND3X1_86 gnd vdd FILL
XFILL_76_DFFSR_192 gnd vdd FILL
XFILL_50_DFFSR_106 gnd vdd FILL
XFILL_27_DFFSR_205 gnd vdd FILL
XFILL_6_BUFX4_31 gnd vdd FILL
XFILL_6_BUFX4_42 gnd vdd FILL
XFILL_6_NAND3X1_97 gnd vdd FILL
XFILL_50_DFFSR_117 gnd vdd FILL
XFILL_27_DFFSR_216 gnd vdd FILL
XFILL_50_DFFSR_128 gnd vdd FILL
XFILL_6_BUFX4_53 gnd vdd FILL
XFILL_27_DFFSR_227 gnd vdd FILL
XFILL_6_BUFX4_64 gnd vdd FILL
XFILL_27_DFFSR_238 gnd vdd FILL
XFILL_41_DFFSR_18 gnd vdd FILL
XFILL_50_DFFSR_139 gnd vdd FILL
XFILL_27_DFFSR_249 gnd vdd FILL
XFILL_41_DFFSR_29 gnd vdd FILL
XFILL_6_BUFX4_75 gnd vdd FILL
XFILL_6_BUFX4_86 gnd vdd FILL
XFILL_6_BUFX4_97 gnd vdd FILL
XFILL_54_DFFSR_105 gnd vdd FILL
XFILL_18_CLKBUF1_19 gnd vdd FILL
XFILL_8_BUFX2_5 gnd vdd FILL
XFILL_54_DFFSR_116 gnd vdd FILL
XFILL_54_DFFSR_127 gnd vdd FILL
XFILL_54_DFFSR_138 gnd vdd FILL
XFILL_81_DFFSR_17 gnd vdd FILL
XFILL_54_DFFSR_149 gnd vdd FILL
XFILL_13_AOI21X1_16 gnd vdd FILL
XFILL_81_DFFSR_28 gnd vdd FILL
XFILL_81_DFFSR_39 gnd vdd FILL
XFILL_13_AOI21X1_27 gnd vdd FILL
XFILL_13_AOI21X1_38 gnd vdd FILL
XFILL_13_AOI21X1_49 gnd vdd FILL
XFILL_10_DFFSR_17 gnd vdd FILL
XFILL_58_DFFSR_104 gnd vdd FILL
XFILL_10_DFFSR_28 gnd vdd FILL
XFILL_10_DFFSR_39 gnd vdd FILL
XFILL_58_DFFSR_115 gnd vdd FILL
XFILL_58_DFFSR_126 gnd vdd FILL
XFILL_58_DFFSR_137 gnd vdd FILL
XFILL_67_DFFSR_4 gnd vdd FILL
XFILL_58_DFFSR_148 gnd vdd FILL
XFILL_58_DFFSR_159 gnd vdd FILL
XFILL_6_OR2X2_1 gnd vdd FILL
XFILL_1_DFFSR_108 gnd vdd FILL
XFILL_50_DFFSR_16 gnd vdd FILL
XFILL_50_DFFSR_27 gnd vdd FILL
XFILL_1_DFFSR_119 gnd vdd FILL
XFILL_50_DFFSR_38 gnd vdd FILL
XFILL_8_5_1 gnd vdd FILL
XFILL_50_DFFSR_49 gnd vdd FILL
XFILL_7_0_0 gnd vdd FILL
XFILL_12_DFFSR_260 gnd vdd FILL
XFILL_5_DFFSR_107 gnd vdd FILL
XFILL_12_DFFSR_271 gnd vdd FILL
XFILL_7_MUX2X1_8 gnd vdd FILL
XFILL_5_DFFSR_118 gnd vdd FILL
XFILL_25_CLKBUF1_10 gnd vdd FILL
XFILL_5_DFFSR_129 gnd vdd FILL
XFILL_25_CLKBUF1_21 gnd vdd FILL
XFILL_25_CLKBUF1_32 gnd vdd FILL
XFILL_0_AOI21X1_3 gnd vdd FILL
XFILL_10_BUFX4_80 gnd vdd FILL
XFILL_16_DFFSR_270 gnd vdd FILL
XFILL_8_CLKBUF1_14 gnd vdd FILL
XFILL_9_DFFSR_106 gnd vdd FILL
XFILL_10_BUFX4_91 gnd vdd FILL
XFILL_8_CLKBUF1_25 gnd vdd FILL
XFILL_9_DFFSR_117 gnd vdd FILL
XFILL_13_MUX2X1_15 gnd vdd FILL
XFILL_8_CLKBUF1_36 gnd vdd FILL
XFILL_9_DFFSR_128 gnd vdd FILL
XFILL_13_MUX2X1_26 gnd vdd FILL
XFILL_3_AOI21X1_11 gnd vdd FILL
XFILL_13_MUX2X1_37 gnd vdd FILL
XFILL_16_4_1 gnd vdd FILL
XFILL_9_DFFSR_139 gnd vdd FILL
XFILL_4_AOI21X1_2 gnd vdd FILL
XFILL_3_AOI21X1_22 gnd vdd FILL
XFILL_13_MUX2X1_48 gnd vdd FILL
XFILL_3_AOI21X1_33 gnd vdd FILL
XFILL_13_MUX2X1_59 gnd vdd FILL
XFILL_3_AOI21X1_44 gnd vdd FILL
XFILL_3_AOI21X1_55 gnd vdd FILL
XFILL_43_DFFSR_170 gnd vdd FILL
XOAI21X1_14 MUX2X1_90/B OAI21X1_4/B OAI21X1_14/C gnd NOR2X1_76/A vdd OAI21X1
XFILL_3_AOI21X1_66 gnd vdd FILL
XFILL_1_NOR3X1_19 gnd vdd FILL
XFILL_13_OAI22X1_13 gnd vdd FILL
XOAI21X1_25 INVX1_194/Y OAI21X1_6/B OAI21X1_25/C gnd NOR2X1_95/B vdd OAI21X1
XFILL_13_OAI22X1_24 gnd vdd FILL
XFILL_43_DFFSR_181 gnd vdd FILL
XFILL_13_OAI22X1_35 gnd vdd FILL
XFILL_3_AOI21X1_77 gnd vdd FILL
XFILL_17_MUX2X1_14 gnd vdd FILL
XFILL_43_DFFSR_192 gnd vdd FILL
XFILL_17_MUX2X1_25 gnd vdd FILL
XFILL_13_OAI22X1_46 gnd vdd FILL
XOAI21X1_36 OAI21X1_1/A OAI21X1_1/B AND2X2_8/B gnd OAI21X1_36/Y vdd OAI21X1
XFILL_17_MUX2X1_36 gnd vdd FILL
XOAI21X1_47 OAI21X1_47/A NOR3X1_48/Y NOR3X1_9/A gnd NOR2X1_44/B vdd OAI21X1
XFILL_17_MUX2X1_47 gnd vdd FILL
XFILL_6_NOR2X1_110 gnd vdd FILL
XFILL_8_AOI21X1_1 gnd vdd FILL
XFILL_6_NOR2X1_121 gnd vdd FILL
XFILL_6_NOR2X1_132 gnd vdd FILL
XFILL_17_MUX2X1_58 gnd vdd FILL
XFILL_17_MUX2X1_69 gnd vdd FILL
XFILL_13_NAND3X1_101 gnd vdd FILL
XFILL_6_NOR2X1_143 gnd vdd FILL
XFILL_2_DFFSR_16 gnd vdd FILL
XFILL_5_NOR3X1_18 gnd vdd FILL
XFILL_2_DFFSR_27 gnd vdd FILL
XFILL_6_NOR2X1_154 gnd vdd FILL
XFILL_13_NAND3X1_112 gnd vdd FILL
XFILL_2_DFFSR_38 gnd vdd FILL
XFILL_47_DFFSR_180 gnd vdd FILL
XFILL_6_NOR2X1_165 gnd vdd FILL
XFILL_2_DFFSR_49 gnd vdd FILL
XFILL_13_NAND3X1_123 gnd vdd FILL
XFILL_5_NOR3X1_29 gnd vdd FILL
XFILL_6_INVX1_3 gnd vdd FILL
XFILL_6_NOR2X1_176 gnd vdd FILL
XFILL_47_DFFSR_191 gnd vdd FILL
XFILL_6_NOR2X1_187 gnd vdd FILL
XFILL_21_DFFSR_105 gnd vdd FILL
XFILL_6_NOR2X1_198 gnd vdd FILL
XFILL_21_DFFSR_116 gnd vdd FILL
XFILL_21_DFFSR_127 gnd vdd FILL
XFILL_21_DFFSR_138 gnd vdd FILL
XFILL_4_INVX1_70 gnd vdd FILL
XFILL_10_NOR2X1_204 gnd vdd FILL
XFILL_21_DFFSR_149 gnd vdd FILL
XFILL_9_NOR3X1_17 gnd vdd FILL
XFILL_4_INVX1_81 gnd vdd FILL
XFILL_4_INVX1_92 gnd vdd FILL
XFILL_9_NOR3X1_28 gnd vdd FILL
XFILL_9_NOR3X1_39 gnd vdd FILL
XFILL_25_DFFSR_104 gnd vdd FILL
XFILL_11_MUX2X1_2 gnd vdd FILL
XFILL_25_DFFSR_115 gnd vdd FILL
XFILL_25_DFFSR_126 gnd vdd FILL
XFILL_23_MUX2X1_101 gnd vdd FILL
XFILL_25_DFFSR_137 gnd vdd FILL
XFILL_23_MUX2X1_112 gnd vdd FILL
XFILL_23_MUX2X1_123 gnd vdd FILL
XFILL_25_DFFSR_148 gnd vdd FILL
XFILL_23_MUX2X1_134 gnd vdd FILL
XFILL_23_MUX2X1_145 gnd vdd FILL
XFILL_25_DFFSR_159 gnd vdd FILL
XFILL_4_NAND3X1_106 gnd vdd FILL
XFILL_4_NAND3X1_117 gnd vdd FILL
XFILL_4_NAND3X1_128 gnd vdd FILL
XFILL_23_MUX2X1_156 gnd vdd FILL
XFILL_29_DFFSR_103 gnd vdd FILL
XFILL_23_MUX2X1_167 gnd vdd FILL
XFILL_6_MUX2X1_105 gnd vdd FILL
XFILL_6_MUX2X1_116 gnd vdd FILL
XFILL_23_MUX2X1_178 gnd vdd FILL
XFILL_23_MUX2X1_189 gnd vdd FILL
XFILL_29_DFFSR_114 gnd vdd FILL
XFILL_6_MUX2X1_127 gnd vdd FILL
XFILL_29_DFFSR_125 gnd vdd FILL
XFILL_29_DFFSR_136 gnd vdd FILL
XFILL_6_MUX2X1_138 gnd vdd FILL
XFILL_6_MUX2X1_149 gnd vdd FILL
XFILL_29_DFFSR_147 gnd vdd FILL
XFILL_19_DFFSR_50 gnd vdd FILL
XFILL_2_BUFX4_90 gnd vdd FILL
XFILL_29_DFFSR_158 gnd vdd FILL
XFILL_19_DFFSR_61 gnd vdd FILL
XFILL_66_3_1 gnd vdd FILL
XFILL_3_OAI22X1_30 gnd vdd FILL
XFILL_29_DFFSR_169 gnd vdd FILL
XFILL_19_DFFSR_72 gnd vdd FILL
XFILL_19_DFFSR_83 gnd vdd FILL
XFILL_21_NOR3X1_16 gnd vdd FILL
XFILL_3_OAI22X1_41 gnd vdd FILL
XFILL_19_DFFSR_94 gnd vdd FILL
XFILL_21_NOR3X1_27 gnd vdd FILL
XFILL_7_OAI21X1_10 gnd vdd FILL
XFILL_7_OAI21X1_21 gnd vdd FILL
XFILL_21_NOR3X1_38 gnd vdd FILL
XFILL_21_NOR3X1_49 gnd vdd FILL
XFILL_71_DFFSR_205 gnd vdd FILL
XFILL_7_OAI21X1_32 gnd vdd FILL
XFILL_7_OAI21X1_43 gnd vdd FILL
XFILL_71_DFFSR_216 gnd vdd FILL
XFILL_71_DFFSR_227 gnd vdd FILL
XFILL_59_DFFSR_60 gnd vdd FILL
XFILL_71_DFFSR_238 gnd vdd FILL
XFILL_71_DFFSR_249 gnd vdd FILL
XFILL_59_DFFSR_71 gnd vdd FILL
XFILL_59_DFFSR_82 gnd vdd FILL
XFILL_25_NOR3X1_15 gnd vdd FILL
XFILL_59_DFFSR_93 gnd vdd FILL
XFILL_25_NOR3X1_26 gnd vdd FILL
XFILL_25_NOR3X1_37 gnd vdd FILL
XFILL_25_NOR3X1_48 gnd vdd FILL
XFILL_75_DFFSR_204 gnd vdd FILL
XFILL_4_NOR2X1_3 gnd vdd FILL
XFILL_75_DFFSR_215 gnd vdd FILL
XFILL_50_7_2 gnd vdd FILL
XFILL_75_DFFSR_226 gnd vdd FILL
XFILL_75_DFFSR_237 gnd vdd FILL
XFILL_75_DFFSR_248 gnd vdd FILL
XFILL_10_DFFSR_170 gnd vdd FILL
XFILL_29_NOR3X1_14 gnd vdd FILL
XFILL_75_DFFSR_259 gnd vdd FILL
XFILL_29_NOR3X1_25 gnd vdd FILL
XFILL_10_DFFSR_181 gnd vdd FILL
XFILL_10_DFFSR_192 gnd vdd FILL
XFILL_29_NOR3X1_36 gnd vdd FILL
XFILL_28_DFFSR_70 gnd vdd FILL
XFILL_29_NOR3X1_47 gnd vdd FILL
XFILL_79_DFFSR_203 gnd vdd FILL
XFILL_28_DFFSR_81 gnd vdd FILL
XFILL_79_DFFSR_214 gnd vdd FILL
XFILL_28_DFFSR_92 gnd vdd FILL
XFILL_79_DFFSR_225 gnd vdd FILL
XFILL_79_DFFSR_236 gnd vdd FILL
XFILL_79_DFFSR_247 gnd vdd FILL
XFILL_3_MUX2X1_1 gnd vdd FILL
XFILL_3_CLKBUF1_1 gnd vdd FILL
XFILL_79_DFFSR_258 gnd vdd FILL
XFILL_14_DFFSR_180 gnd vdd FILL
XFILL_79_DFFSR_269 gnd vdd FILL
XFILL_14_DFFSR_191 gnd vdd FILL
XFILL_68_DFFSR_80 gnd vdd FILL
XFILL_11_DFFSR_3 gnd vdd FILL
XFILL_9_NAND3X1_19 gnd vdd FILL
XFILL_68_DFFSR_91 gnd vdd FILL
XFILL_49_DFFSR_1 gnd vdd FILL
XFILL_18_DFFSR_190 gnd vdd FILL
XFILL_0_NOR3X1_7 gnd vdd FILL
XFILL_37_DFFSR_90 gnd vdd FILL
XFILL_60_DFFSR_270 gnd vdd FILL
XFILL_57_3_1 gnd vdd FILL
XFILL_33_DFFSR_7 gnd vdd FILL
XFILL_0_OAI21X1_6 gnd vdd FILL
XFILL_12_MUX2X1_130 gnd vdd FILL
XFILL_12_MUX2X1_141 gnd vdd FILL
XFILL_12_MUX2X1_152 gnd vdd FILL
XFILL_12_MUX2X1_163 gnd vdd FILL
XFILL_41_7_2 gnd vdd FILL
XFILL_12_MUX2X1_174 gnd vdd FILL
XFILL_12_MUX2X1_185 gnd vdd FILL
XFILL_42_DFFSR_204 gnd vdd FILL
XFILL_40_2_1 gnd vdd FILL
XFILL_42_DFFSR_215 gnd vdd FILL
XFILL_4_OAI21X1_5 gnd vdd FILL
XFILL_1_NOR2X1_30 gnd vdd FILL
XFILL_1_NOR2X1_41 gnd vdd FILL
XFILL_42_DFFSR_226 gnd vdd FILL
XFILL_1_NOR2X1_52 gnd vdd FILL
XFILL_42_DFFSR_237 gnd vdd FILL
XFILL_42_DFFSR_248 gnd vdd FILL
XFILL_1_NOR2X1_63 gnd vdd FILL
XFILL_42_DFFSR_259 gnd vdd FILL
XFILL_1_NOR2X1_74 gnd vdd FILL
XFILL_1_NOR2X1_85 gnd vdd FILL
XFILL_1_NOR2X1_96 gnd vdd FILL
XFILL_46_DFFSR_203 gnd vdd FILL
XFILL_46_DFFSR_214 gnd vdd FILL
XFILL_8_OAI21X1_4 gnd vdd FILL
XFILL_46_DFFSR_225 gnd vdd FILL
XFILL_5_NOR2X1_40 gnd vdd FILL
XFILL_5_NOR2X1_51 gnd vdd FILL
XFILL_46_DFFSR_236 gnd vdd FILL
XFILL_5_NOR2X1_62 gnd vdd FILL
XFILL_46_DFFSR_247 gnd vdd FILL
XFILL_46_DFFSR_258 gnd vdd FILL
XFILL_46_DFFSR_269 gnd vdd FILL
XFILL_5_NOR2X1_73 gnd vdd FILL
XFILL_5_NOR2X1_84 gnd vdd FILL
XFILL_5_NOR2X1_95 gnd vdd FILL
XFILL_73_DFFSR_103 gnd vdd FILL
XFILL_73_DFFSR_114 gnd vdd FILL
XFILL_73_DFFSR_125 gnd vdd FILL
XFILL_73_DFFSR_136 gnd vdd FILL
XFILL_13_OAI22X1_1 gnd vdd FILL
XFILL_73_DFFSR_147 gnd vdd FILL
XFILL_9_NOR2X1_50 gnd vdd FILL
XFILL_9_NOR2X1_61 gnd vdd FILL
XFILL_73_DFFSR_158 gnd vdd FILL
XFILL_73_DFFSR_169 gnd vdd FILL
XFILL_9_NOR2X1_72 gnd vdd FILL
XFILL_9_NOR2X1_83 gnd vdd FILL
XFILL_77_DFFSR_102 gnd vdd FILL
XFILL_9_NOR2X1_94 gnd vdd FILL
XFILL_6_7 gnd vdd FILL
XFILL_77_DFFSR_113 gnd vdd FILL
XFILL_77_DFFSR_124 gnd vdd FILL
XFILL_9_NOR2X1_109 gnd vdd FILL
XFILL_77_DFFSR_135 gnd vdd FILL
XFILL_77_DFFSR_146 gnd vdd FILL
XFILL_15_NAND3X1_11 gnd vdd FILL
XFILL_77_DFFSR_157 gnd vdd FILL
XFILL_15_NAND3X1_22 gnd vdd FILL
XFILL_48_3_1 gnd vdd FILL
XFILL_77_DFFSR_168 gnd vdd FILL
XFILL_15_NAND3X1_33 gnd vdd FILL
XFILL_2_MUX2X1_180 gnd vdd FILL
XFILL_77_DFFSR_179 gnd vdd FILL
XFILL_15_NAND3X1_44 gnd vdd FILL
XFILL_2_MUX2X1_191 gnd vdd FILL
XFILL_15_NAND3X1_55 gnd vdd FILL
XFILL_15_NAND3X1_66 gnd vdd FILL
XFILL_35_CLKBUF1_11 gnd vdd FILL
XFILL_35_CLKBUF1_22 gnd vdd FILL
XFILL_15_NAND3X1_77 gnd vdd FILL
XFILL_14_AND2X2_8 gnd vdd FILL
XFILL_15_NAND3X1_88 gnd vdd FILL
XFILL_35_CLKBUF1_33 gnd vdd FILL
XFILL_15_NAND3X1_99 gnd vdd FILL
XFILL_1_NAND2X1_7 gnd vdd FILL
XFILL_32_7_2 gnd vdd FILL
XFILL_11_BUFX4_14 gnd vdd FILL
XFILL_11_BUFX4_25 gnd vdd FILL
XFILL_31_2_1 gnd vdd FILL
XFILL_11_BUFX4_36 gnd vdd FILL
XFILL_11_BUFX4_47 gnd vdd FILL
XFILL_5_NAND2X1_6 gnd vdd FILL
XFILL_11_BUFX4_58 gnd vdd FILL
XFILL_11_BUFX4_69 gnd vdd FILL
XFILL_6_OAI22X1_18 gnd vdd FILL
XFILL_1_MUX2X1_70 gnd vdd FILL
XFILL_1_MUX2X1_81 gnd vdd FILL
XFILL_14_NAND3X1_102 gnd vdd FILL
XFILL_1_MUX2X1_92 gnd vdd FILL
XFILL_14_NAND3X1_113 gnd vdd FILL
XFILL_6_OAI22X1_29 gnd vdd FILL
XDFFSR_17 DFFSR_17/Q DFFSR_88/CLK DFFSR_87/R vdd DFFSR_17/D gnd vdd DFFSR
XFILL_14_NAND3X1_124 gnd vdd FILL
XFILL_62_DFFSR_190 gnd vdd FILL
XDFFSR_28 DFFSR_28/Q DFFSR_4/CLK DFFSR_4/R vdd DFFSR_28/D gnd vdd DFFSR
XFILL_9_NAND2X1_5 gnd vdd FILL
XFILL_19_AOI22X1_11 gnd vdd FILL
XDFFSR_39 INVX1_23/A DFFSR_39/CLK DFFSR_45/R vdd DFFSR_39/D gnd vdd DFFSR
XFILL_13_DFFSR_203 gnd vdd FILL
XFILL_10_NAND3X1_3 gnd vdd FILL
XFILL_13_DFFSR_214 gnd vdd FILL
XFILL_13_DFFSR_225 gnd vdd FILL
XFILL_13_DFFSR_236 gnd vdd FILL
XFILL_5_MUX2X1_80 gnd vdd FILL
XFILL_13_DFFSR_247 gnd vdd FILL
XFILL_5_MUX2X1_91 gnd vdd FILL
XFILL_5_NAND3X1_50 gnd vdd FILL
XFILL_13_DFFSR_258 gnd vdd FILL
XFILL_50_DFFSR_1 gnd vdd FILL
XFILL_5_NAND3X1_61 gnd vdd FILL
XFILL_13_DFFSR_269 gnd vdd FILL
XFILL_5_NAND3X1_72 gnd vdd FILL
XFILL_5_NAND3X1_83 gnd vdd FILL
XFILL_9_NAND2X1_30 gnd vdd FILL
XFILL_17_DFFSR_202 gnd vdd FILL
XFILL_5_NAND3X1_94 gnd vdd FILL
XFILL_40_DFFSR_103 gnd vdd FILL
XFILL_9_NAND2X1_41 gnd vdd FILL
XFILL_17_DFFSR_213 gnd vdd FILL
XFILL_9_NAND2X1_52 gnd vdd FILL
XFILL_40_DFFSR_114 gnd vdd FILL
XFILL_14_NAND3X1_2 gnd vdd FILL
XFILL_9_NAND2X1_63 gnd vdd FILL
XFILL_40_DFFSR_125 gnd vdd FILL
XFILL_40_DFFSR_136 gnd vdd FILL
XFILL_9_NAND2X1_74 gnd vdd FILL
XFILL_17_DFFSR_224 gnd vdd FILL
XFILL_17_DFFSR_235 gnd vdd FILL
XFILL_5_INVX1_15 gnd vdd FILL
XFILL_5_NAND3X1_107 gnd vdd FILL
XFILL_5_INVX1_26 gnd vdd FILL
XFILL_9_NAND2X1_85 gnd vdd FILL
XCLKBUF1_15 BUFX4_84/Y gnd DFFSR_78/CLK vdd CLKBUF1
XFILL_22_12 gnd vdd FILL
XFILL_17_DFFSR_246 gnd vdd FILL
XFILL_40_DFFSR_147 gnd vdd FILL
XFILL_40_DFFSR_158 gnd vdd FILL
XFILL_5_INVX1_37 gnd vdd FILL
XFILL_9_MUX2X1_90 gnd vdd FILL
XFILL_9_NAND2X1_96 gnd vdd FILL
XFILL_17_DFFSR_257 gnd vdd FILL
XFILL_17_DFFSR_268 gnd vdd FILL
XFILL_5_NAND3X1_118 gnd vdd FILL
XFILL_5_INVX1_48 gnd vdd FILL
XFILL_40_DFFSR_169 gnd vdd FILL
XCLKBUF1_26 BUFX4_4/Y gnd CLKBUF1_26/Y vdd CLKBUF1
XFILL_5_NAND3X1_129 gnd vdd FILL
XFILL_6_AND2X2_7 gnd vdd FILL
XCLKBUF1_37 BUFX4_9/Y gnd DFFSR_39/CLK vdd CLKBUF1
XFILL_5_INVX1_59 gnd vdd FILL
XFILL_44_DFFSR_102 gnd vdd FILL
XFILL_17_CLKBUF1_16 gnd vdd FILL
XFILL_44_DFFSR_113 gnd vdd FILL
XFILL_44_DFFSR_124 gnd vdd FILL
XFILL_39_3_1 gnd vdd FILL
XFILL_17_CLKBUF1_27 gnd vdd FILL
XFILL_17_CLKBUF1_38 gnd vdd FILL
XFILL_44_DFFSR_135 gnd vdd FILL
XFILL_44_DFFSR_146 gnd vdd FILL
XFILL_12_AOI21X1_13 gnd vdd FILL
XFILL_44_DFFSR_157 gnd vdd FILL
XFILL_12_AOI21X1_24 gnd vdd FILL
XBUFX4_80 INVX8_4/Y gnd BUFX4_80/Y vdd BUFX4
XFILL_44_DFFSR_168 gnd vdd FILL
XFILL_12_AOI21X1_35 gnd vdd FILL
XFILL_12_AOI21X1_46 gnd vdd FILL
XFILL_44_DFFSR_179 gnd vdd FILL
XBUFX4_91 BUFX4_92/A gnd BUFX4_91/Y vdd BUFX4
XFILL_48_DFFSR_101 gnd vdd FILL
XFILL_2_DFFSR_6 gnd vdd FILL
XFILL_12_AOI21X1_57 gnd vdd FILL
XFILL_15_DFFSR_4 gnd vdd FILL
XFILL_12_AOI21X1_68 gnd vdd FILL
XFILL_48_DFFSR_112 gnd vdd FILL
XFILL_3_BUFX4_13 gnd vdd FILL
XFILL_12_AOI21X1_79 gnd vdd FILL
XFILL_48_DFFSR_123 gnd vdd FILL
XFILL_72_DFFSR_5 gnd vdd FILL
XFILL_48_DFFSR_134 gnd vdd FILL
XFILL_3_BUFX4_24 gnd vdd FILL
XFILL_48_DFFSR_145 gnd vdd FILL
XFILL_3_BUFX4_35 gnd vdd FILL
XFILL_48_DFFSR_156 gnd vdd FILL
XFILL_3_BUFX4_46 gnd vdd FILL
XFILL_10_AOI22X1_8 gnd vdd FILL
XFILL_3_BUFX4_57 gnd vdd FILL
XFILL_48_DFFSR_167 gnd vdd FILL
XFILL_3_BUFX4_68 gnd vdd FILL
XFILL_48_DFFSR_178 gnd vdd FILL
XFILL_48_DFFSR_189 gnd vdd FILL
XFILL_3_BUFX4_79 gnd vdd FILL
XFILL_23_7_2 gnd vdd FILL
XFILL_22_2_1 gnd vdd FILL
XFILL_14_AOI22X1_7 gnd vdd FILL
XFILL_0_NAND3X1_103 gnd vdd FILL
XFILL_24_CLKBUF1_40 gnd vdd FILL
XFILL_18_AOI22X1_6 gnd vdd FILL
XFILL_0_NAND3X1_114 gnd vdd FILL
XFILL_0_NAND3X1_125 gnd vdd FILL
XFILL_7_CLKBUF1_11 gnd vdd FILL
XFILL_37_DFFSR_8 gnd vdd FILL
XFILL_7_CLKBUF1_22 gnd vdd FILL
XFILL_10_AND2X2_1 gnd vdd FILL
XFILL_7_CLKBUF1_33 gnd vdd FILL
XFILL_29_DFFSR_15 gnd vdd FILL
XFILL_29_DFFSR_26 gnd vdd FILL
XFILL_29_DFFSR_37 gnd vdd FILL
XFILL_15_MUX2X1_107 gnd vdd FILL
XFILL_15_MUX2X1_118 gnd vdd FILL
XFILL_29_DFFSR_48 gnd vdd FILL
XFILL_15_MUX2X1_129 gnd vdd FILL
XFILL_2_AOI21X1_30 gnd vdd FILL
XFILL_29_DFFSR_59 gnd vdd FILL
XFILL_2_AOI21X1_41 gnd vdd FILL
XFILL_2_AOI21X1_52 gnd vdd FILL
XFILL_12_OAI22X1_10 gnd vdd FILL
XFILL_2_AOI21X1_63 gnd vdd FILL
XFILL_12_OAI22X1_21 gnd vdd FILL
XFILL_2_AOI21X1_74 gnd vdd FILL
XFILL_69_DFFSR_14 gnd vdd FILL
XFILL_12_OAI22X1_32 gnd vdd FILL
XFILL_12_OAI22X1_43 gnd vdd FILL
XFILL_69_DFFSR_25 gnd vdd FILL
XFILL_69_DFFSR_36 gnd vdd FILL
XFILL_69_DFFSR_47 gnd vdd FILL
XFILL_69_DFFSR_58 gnd vdd FILL
XFILL_69_DFFSR_69 gnd vdd FILL
XFILL_5_NOR2X1_140 gnd vdd FILL
XFILL_5_NOR2X1_151 gnd vdd FILL
XFILL_5_NOR2X1_162 gnd vdd FILL
XFILL_5_3_1 gnd vdd FILL
XFILL_5_NOR2X1_173 gnd vdd FILL
XFILL_11_DFFSR_102 gnd vdd FILL
XFILL_5_NOR2X1_184 gnd vdd FILL
XFILL_5_NOR2X1_195 gnd vdd FILL
XFILL_11_DFFSR_113 gnd vdd FILL
XFILL_11_DFFSR_124 gnd vdd FILL
XFILL_11_DFFSR_135 gnd vdd FILL
XFILL_38_DFFSR_13 gnd vdd FILL
XFILL_11_DFFSR_146 gnd vdd FILL
XFILL_38_DFFSR_24 gnd vdd FILL
XFILL_11_DFFSR_157 gnd vdd FILL
XFILL_38_DFFSR_35 gnd vdd FILL
XFILL_11_DFFSR_168 gnd vdd FILL
XFILL_11_DFFSR_179 gnd vdd FILL
XFILL_38_DFFSR_46 gnd vdd FILL
XFILL_15_DFFSR_101 gnd vdd FILL
XFILL_38_DFFSR_57 gnd vdd FILL
XFILL_38_DFFSR_68 gnd vdd FILL
XFILL_38_DFFSR_79 gnd vdd FILL
XFILL_15_DFFSR_112 gnd vdd FILL
XFILL_15_DFFSR_123 gnd vdd FILL
XFILL_15_DFFSR_134 gnd vdd FILL
XFILL_22_MUX2X1_120 gnd vdd FILL
XFILL_78_DFFSR_12 gnd vdd FILL
XFILL_15_DFFSR_145 gnd vdd FILL
XFILL_14_7_2 gnd vdd FILL
XFILL_22_MUX2X1_131 gnd vdd FILL
XFILL_78_DFFSR_23 gnd vdd FILL
XFILL_15_DFFSR_156 gnd vdd FILL
XFILL_22_MUX2X1_142 gnd vdd FILL
XFILL_78_DFFSR_34 gnd vdd FILL
XFILL_22_MUX2X1_153 gnd vdd FILL
XFILL_15_DFFSR_167 gnd vdd FILL
XFILL_15_DFFSR_178 gnd vdd FILL
XFILL_13_2_1 gnd vdd FILL
XFILL_78_DFFSR_45 gnd vdd FILL
XFILL_78_DFFSR_56 gnd vdd FILL
XFILL_5_MUX2X1_102 gnd vdd FILL
XFILL_22_MUX2X1_164 gnd vdd FILL
XFILL_19_DFFSR_100 gnd vdd FILL
XFILL_15_DFFSR_189 gnd vdd FILL
XFILL_22_MUX2X1_175 gnd vdd FILL
XFILL_5_MUX2X1_113 gnd vdd FILL
XFILL_78_DFFSR_67 gnd vdd FILL
XFILL_5_MUX2X1_124 gnd vdd FILL
XFILL_78_DFFSR_78 gnd vdd FILL
XFILL_22_MUX2X1_186 gnd vdd FILL
XFILL_19_DFFSR_111 gnd vdd FILL
XFILL_78_DFFSR_89 gnd vdd FILL
XFILL_19_DFFSR_122 gnd vdd FILL
XFILL_19_DFFSR_133 gnd vdd FILL
XFILL_5_MUX2X1_135 gnd vdd FILL
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XFILL_5_MUX2X1_146 gnd vdd FILL
XFILL_19_DFFSR_144 gnd vdd FILL
XFILL_1_INVX1_30 gnd vdd FILL
XFILL_19_DFFSR_155 gnd vdd FILL
XFILL_1_INVX1_41 gnd vdd FILL
XFILL_5_MUX2X1_157 gnd vdd FILL
XFILL_1_INVX1_52 gnd vdd FILL
XFILL_5_MUX2X1_168 gnd vdd FILL
XFILL_0_BUFX4_105 gnd vdd FILL
XFILL_19_DFFSR_166 gnd vdd FILL
XFILL_1_INVX1_63 gnd vdd FILL
XFILL_8_CLKBUF1_9 gnd vdd FILL
XFILL_19_DFFSR_177 gnd vdd FILL
XFILL_11_NOR3X1_13 gnd vdd FILL
XFILL_1_INVX1_74 gnd vdd FILL
XFILL_5_MUX2X1_179 gnd vdd FILL
XFILL_47_DFFSR_11 gnd vdd FILL
XFILL_11_NOR3X1_24 gnd vdd FILL
XFILL_19_DFFSR_188 gnd vdd FILL
XFILL_1_INVX1_85 gnd vdd FILL
XFILL_47_DFFSR_22 gnd vdd FILL
XFILL_19_DFFSR_199 gnd vdd FILL
XFILL_1_INVX1_96 gnd vdd FILL
XFILL_11_NOR3X1_35 gnd vdd FILL
XFILL_47_DFFSR_33 gnd vdd FILL
XFILL_61_DFFSR_202 gnd vdd FILL
XFILL_18_NOR3X1_8 gnd vdd FILL
XFILL_11_NOR3X1_46 gnd vdd FILL
XFILL_47_DFFSR_44 gnd vdd FILL
XFILL_61_DFFSR_213 gnd vdd FILL
XFILL_6_OAI21X1_40 gnd vdd FILL
XFILL_47_DFFSR_55 gnd vdd FILL
XFILL_4_BUFX4_104 gnd vdd FILL
XFILL_47_DFFSR_66 gnd vdd FILL
XFILL_61_DFFSR_224 gnd vdd FILL
XFILL_47_DFFSR_77 gnd vdd FILL
XFILL_61_DFFSR_235 gnd vdd FILL
XFILL_47_DFFSR_88 gnd vdd FILL
XFILL_61_DFFSR_246 gnd vdd FILL
XFILL_47_DFFSR_99 gnd vdd FILL
XFILL_15_NOR3X1_12 gnd vdd FILL
XFILL_61_DFFSR_257 gnd vdd FILL
XFILL_15_NOR3X1_23 gnd vdd FILL
XFILL_87_DFFSR_10 gnd vdd FILL
XFILL_61_DFFSR_268 gnd vdd FILL
XFILL_87_DFFSR_21 gnd vdd FILL
XFILL_15_NOR3X1_34 gnd vdd FILL
XFILL_87_DFFSR_32 gnd vdd FILL
XFILL_65_DFFSR_201 gnd vdd FILL
XFILL_87_DFFSR_43 gnd vdd FILL
XFILL_15_NOR3X1_45 gnd vdd FILL
XFILL_65_DFFSR_212 gnd vdd FILL
XFILL_87_DFFSR_54 gnd vdd FILL
XFILL_65_DFFSR_223 gnd vdd FILL
XFILL_16_DFFSR_10 gnd vdd FILL
XFILL_16_DFFSR_21 gnd vdd FILL
XFILL_87_DFFSR_65 gnd vdd FILL
XFILL_8_BUFX4_103 gnd vdd FILL
XFILL_87_DFFSR_76 gnd vdd FILL
XFILL_65_DFFSR_234 gnd vdd FILL
XFILL_16_DFFSR_32 gnd vdd FILL
XFILL_16_DFFSR_43 gnd vdd FILL
XFILL_87_DFFSR_87 gnd vdd FILL
XFILL_65_DFFSR_245 gnd vdd FILL
XFILL_19_NOR3X1_11 gnd vdd FILL
XFILL_87_DFFSR_98 gnd vdd FILL
XFILL_4_4 gnd vdd FILL
XFILL_65_DFFSR_256 gnd vdd FILL
XFILL_16_DFFSR_54 gnd vdd FILL
XFILL_12_INVX8_2 gnd vdd FILL
XFILL_65_DFFSR_267 gnd vdd FILL
XFILL_19_NOR3X1_22 gnd vdd FILL
XFILL_19_NOR3X1_33 gnd vdd FILL
XFILL_20_CLKBUF1_8 gnd vdd FILL
XFILL_16_DFFSR_65 gnd vdd FILL
XFILL_16_DFFSR_76 gnd vdd FILL
XFILL_69_DFFSR_200 gnd vdd FILL
XFILL_19_NOR3X1_44 gnd vdd FILL
XFILL_16_DFFSR_87 gnd vdd FILL
XFILL_69_DFFSR_211 gnd vdd FILL
XFILL_16_DFFSR_98 gnd vdd FILL
XFILL_60_6 gnd vdd FILL
XFILL_69_DFFSR_222 gnd vdd FILL
XFILL_56_DFFSR_20 gnd vdd FILL
XFILL_69_DFFSR_233 gnd vdd FILL
XFILL_56_DFFSR_31 gnd vdd FILL
XFILL_27_NOR3X1_6 gnd vdd FILL
XFILL_56_DFFSR_42 gnd vdd FILL
XFILL_69_DFFSR_244 gnd vdd FILL
XFILL_53_5 gnd vdd FILL
XFILL_69_DFFSR_255 gnd vdd FILL
XFILL_56_DFFSR_53 gnd vdd FILL
XFILL_56_DFFSR_64 gnd vdd FILL
XFILL_69_DFFSR_266 gnd vdd FILL
XFILL_24_CLKBUF1_7 gnd vdd FILL
XFILL_64_6_2 gnd vdd FILL
XFILL_56_DFFSR_75 gnd vdd FILL
XFILL_56_DFFSR_86 gnd vdd FILL
XFILL_46_4 gnd vdd FILL
XFILL_56_DFFSR_97 gnd vdd FILL
XFILL_2_NOR2X1_17 gnd vdd FILL
XFILL_63_1_1 gnd vdd FILL
XFILL_8_NAND3X1_16 gnd vdd FILL
XFILL_2_NOR2X1_28 gnd vdd FILL
XFILL_8_NAND3X1_27 gnd vdd FILL
XFILL_2_NOR2X1_39 gnd vdd FILL
XFILL_8_NAND3X1_38 gnd vdd FILL
XFILL_1_NOR2X1_7 gnd vdd FILL
XFILL_54_DFFSR_2 gnd vdd FILL
XFILL_8_NAND3X1_49 gnd vdd FILL
XFILL_28_CLKBUF1_6 gnd vdd FILL
XFILL_25_DFFSR_30 gnd vdd FILL
XFILL_25_DFFSR_41 gnd vdd FILL
XFILL_25_DFFSR_52 gnd vdd FILL
XFILL_6_NOR2X1_16 gnd vdd FILL
XFILL_25_DFFSR_63 gnd vdd FILL
XFILL_6_NOR2X1_27 gnd vdd FILL
XFILL_25_DFFSR_74 gnd vdd FILL
XFILL_6_NOR2X1_38 gnd vdd FILL
XFILL_6_NOR2X1_49 gnd vdd FILL
XFILL_25_DFFSR_85 gnd vdd FILL
XFILL_25_DFFSR_96 gnd vdd FILL
XFILL_65_DFFSR_40 gnd vdd FILL
XFILL_0_MUX2X1_5 gnd vdd FILL
XFILL_65_DFFSR_51 gnd vdd FILL
XFILL_65_DFFSR_62 gnd vdd FILL
XFILL_65_DFFSR_73 gnd vdd FILL
XFILL_65_DFFSR_84 gnd vdd FILL
XFILL_65_DFFSR_95 gnd vdd FILL
XFILL_15_NAND3X1_103 gnd vdd FILL
XFILL_1_NAND2X1_18 gnd vdd FILL
XFILL_15_NAND3X1_114 gnd vdd FILL
XFILL_6_DFFSR_7 gnd vdd FILL
XFILL_1_NAND2X1_29 gnd vdd FILL
XFILL_8_DFFSR_20 gnd vdd FILL
XFILL_15_NAND3X1_125 gnd vdd FILL
XFILL_19_DFFSR_5 gnd vdd FILL
XFILL_8_DFFSR_31 gnd vdd FILL
XFILL_76_DFFSR_6 gnd vdd FILL
XFILL_8_DFFSR_42 gnd vdd FILL
XFILL_8_DFFSR_53 gnd vdd FILL
XFILL_8_DFFSR_64 gnd vdd FILL
XFILL_8_DFFSR_75 gnd vdd FILL
XFILL_18_OAI22X1_9 gnd vdd FILL
XFILL_34_DFFSR_50 gnd vdd FILL
XFILL_8_DFFSR_86 gnd vdd FILL
XFILL_11_MUX2X1_160 gnd vdd FILL
XFILL_34_DFFSR_61 gnd vdd FILL
XFILL_34_DFFSR_72 gnd vdd FILL
XFILL_8_DFFSR_97 gnd vdd FILL
XFILL_34_DFFSR_83 gnd vdd FILL
XFILL_11_MUX2X1_171 gnd vdd FILL
XFILL_34_DFFSR_94 gnd vdd FILL
XFILL_11_MUX2X1_182 gnd vdd FILL
XFILL_32_DFFSR_201 gnd vdd FILL
XFILL_11_MUX2X1_193 gnd vdd FILL
XFILL_32_DFFSR_212 gnd vdd FILL
XFILL_32_DFFSR_223 gnd vdd FILL
XFILL_32_DFFSR_234 gnd vdd FILL
XFILL_6_NAND3X1_108 gnd vdd FILL
XFILL_32_DFFSR_245 gnd vdd FILL
XFILL_74_DFFSR_60 gnd vdd FILL
XFILL_32_DFFSR_256 gnd vdd FILL
XFILL_32_DFFSR_267 gnd vdd FILL
XFILL_6_NAND3X1_119 gnd vdd FILL
XFILL_74_DFFSR_71 gnd vdd FILL
XFILL_74_DFFSR_82 gnd vdd FILL
XFILL_74_DFFSR_93 gnd vdd FILL
XFILL_36_DFFSR_200 gnd vdd FILL
XFILL_36_DFFSR_211 gnd vdd FILL
XFILL_27_CLKBUF1_17 gnd vdd FILL
XFILL_27_CLKBUF1_28 gnd vdd FILL
XFILL_36_DFFSR_222 gnd vdd FILL
XFILL_27_CLKBUF1_39 gnd vdd FILL
XFILL_36_DFFSR_233 gnd vdd FILL
XFILL_55_6_2 gnd vdd FILL
XFILL_36_DFFSR_244 gnd vdd FILL
XFILL_36_DFFSR_255 gnd vdd FILL
XFILL_54_1_1 gnd vdd FILL
XFILL_36_DFFSR_266 gnd vdd FILL
XFILL_2_MUX2X1_13 gnd vdd FILL
XFILL_14_NOR3X1_1 gnd vdd FILL
XFILL_63_DFFSR_100 gnd vdd FILL
XFILL_2_MUX2X1_24 gnd vdd FILL
XFILL_2_MUX2X1_35 gnd vdd FILL
XFILL_63_DFFSR_111 gnd vdd FILL
XFILL_2_MUX2X1_46 gnd vdd FILL
XFILL_5_AOI21X1_18 gnd vdd FILL
XFILL_43_DFFSR_70 gnd vdd FILL
XFILL_2_MUX2X1_57 gnd vdd FILL
XFILL_63_DFFSR_122 gnd vdd FILL
XFILL_63_DFFSR_133 gnd vdd FILL
XFILL_43_DFFSR_81 gnd vdd FILL
XFILL_43_DFFSR_92 gnd vdd FILL
XFILL_63_DFFSR_144 gnd vdd FILL
XFILL_5_AOI21X1_29 gnd vdd FILL
XFILL_2_MUX2X1_68 gnd vdd FILL
XFILL_2_MUX2X1_79 gnd vdd FILL
XFILL_63_DFFSR_155 gnd vdd FILL
XFILL_10_NAND3X1_110 gnd vdd FILL
XFILL_10_NAND3X1_121 gnd vdd FILL
XFILL_63_DFFSR_166 gnd vdd FILL
XFILL_6_MUX2X1_12 gnd vdd FILL
XFILL_63_DFFSR_177 gnd vdd FILL
XFILL_10_NAND3X1_132 gnd vdd FILL
XFILL_6_MUX2X1_23 gnd vdd FILL
XFILL_63_DFFSR_188 gnd vdd FILL
XFILL_6_MUX2X1_34 gnd vdd FILL
XFILL_67_DFFSR_110 gnd vdd FILL
XFILL_63_DFFSR_199 gnd vdd FILL
XFILL_8_NOR2X1_106 gnd vdd FILL
XFILL_6_MUX2X1_45 gnd vdd FILL
XFILL_67_DFFSR_121 gnd vdd FILL
XFILL_6_MUX2X1_56 gnd vdd FILL
XFILL_83_DFFSR_80 gnd vdd FILL
XFILL_67_DFFSR_132 gnd vdd FILL
XFILL_8_NOR2X1_117 gnd vdd FILL
XFILL_67_DFFSR_143 gnd vdd FILL
XFILL_8_NOR2X1_128 gnd vdd FILL
XFILL_83_DFFSR_91 gnd vdd FILL
XFILL_6_MUX2X1_67 gnd vdd FILL
XFILL_67_DFFSR_154 gnd vdd FILL
XFILL_6_MUX2X1_78 gnd vdd FILL
XFILL_8_NOR2X1_139 gnd vdd FILL
XFILL_0_BUFX4_7 gnd vdd FILL
XFILL_14_NAND3X1_30 gnd vdd FILL
XFILL_6_MUX2X1_89 gnd vdd FILL
XFILL_67_DFFSR_165 gnd vdd FILL
XFILL_12_DFFSR_80 gnd vdd FILL
XFILL_14_NAND3X1_41 gnd vdd FILL
XFILL_67_DFFSR_176 gnd vdd FILL
XFILL_13_BUFX4_5 gnd vdd FILL
XFILL_12_DFFSR_91 gnd vdd FILL
XFILL_67_DFFSR_187 gnd vdd FILL
XFILL_14_NAND3X1_52 gnd vdd FILL
XFILL_67_DFFSR_198 gnd vdd FILL
XFILL_14_NAND3X1_63 gnd vdd FILL
XFILL_14_NAND3X1_74 gnd vdd FILL
XFILL_34_CLKBUF1_30 gnd vdd FILL
XFILL_14_NAND3X1_85 gnd vdd FILL
XFILL_34_CLKBUF1_41 gnd vdd FILL
XFILL_14_NAND3X1_96 gnd vdd FILL
XFILL_1_NAND3X1_104 gnd vdd FILL
XFILL_1_NAND3X1_115 gnd vdd FILL
XFILL_1_NAND3X1_126 gnd vdd FILL
XFILL_52_DFFSR_90 gnd vdd FILL
XFILL_11_NOR2X1_90 gnd vdd FILL
XFILL_22_MUX2X1_10 gnd vdd FILL
XFILL_22_MUX2X1_21 gnd vdd FILL
XFILL_22_MUX2X1_32 gnd vdd FILL
XFILL_22_MUX2X1_43 gnd vdd FILL
XFILL_22_MUX2X1_54 gnd vdd FILL
XFILL_5_OAI22X1_15 gnd vdd FILL
XFILL_22_MUX2X1_65 gnd vdd FILL
XFILL_22_MUX2X1_76 gnd vdd FILL
XFILL_5_OAI22X1_26 gnd vdd FILL
XFILL_22_MUX2X1_87 gnd vdd FILL
XFILL_5_OAI22X1_37 gnd vdd FILL
XFILL_22_MUX2X1_98 gnd vdd FILL
XFILL_5_OAI22X1_48 gnd vdd FILL
XFILL_9_OAI21X1_17 gnd vdd FILL
XFILL_46_6_2 gnd vdd FILL
XFILL_9_OAI21X1_28 gnd vdd FILL
XFILL_9_OAI21X1_39 gnd vdd FILL
XFILL_45_1_1 gnd vdd FILL
XFILL_4_NAND3X1_80 gnd vdd FILL
XFILL_4_NAND3X1_91 gnd vdd FILL
XFILL_30_DFFSR_100 gnd vdd FILL
XFILL_30_DFFSR_111 gnd vdd FILL
XFILL_8_NAND2X1_60 gnd vdd FILL
XFILL_2_NOR2X1_206 gnd vdd FILL
XFILL_30_DFFSR_122 gnd vdd FILL
XFILL_30_DFFSR_133 gnd vdd FILL
XFILL_8_NAND2X1_71 gnd vdd FILL
XFILL_4_DFFSR_90 gnd vdd FILL
XFILL_30_DFFSR_144 gnd vdd FILL
XFILL_8_NAND2X1_82 gnd vdd FILL
XFILL_30_DFFSR_155 gnd vdd FILL
XFILL_8_NAND2X1_93 gnd vdd FILL
XFILL_30_DFFSR_166 gnd vdd FILL
XFILL_30_DFFSR_177 gnd vdd FILL
XFILL_16_INVX8_3 gnd vdd FILL
XFILL_30_DFFSR_188 gnd vdd FILL
XFILL_30_DFFSR_199 gnd vdd FILL
XFILL_16_CLKBUF1_13 gnd vdd FILL
XFILL_34_DFFSR_110 gnd vdd FILL
XFILL_11_NAND2X1_1 gnd vdd FILL
XFILL_16_CLKBUF1_24 gnd vdd FILL
XFILL_34_DFFSR_121 gnd vdd FILL
XFILL_34_DFFSR_132 gnd vdd FILL
XFILL_16_CLKBUF1_35 gnd vdd FILL
XFILL_34_DFFSR_143 gnd vdd FILL
XFILL_34_DFFSR_154 gnd vdd FILL
XFILL_11_AOI21X1_10 gnd vdd FILL
XFILL_11_AOI21X1_21 gnd vdd FILL
XFILL_11_AOI21X1_32 gnd vdd FILL
XFILL_34_DFFSR_165 gnd vdd FILL
XFILL_11_AOI21X1_43 gnd vdd FILL
XFILL_34_DFFSR_176 gnd vdd FILL
XAND2X2_1 AND2X2_6/A AND2X2_1/B gnd AND2X2_1/Y vdd AND2X2
XFILL_34_DFFSR_187 gnd vdd FILL
XFILL_11_AOI21X1_54 gnd vdd FILL
XFILL_20_DFFSR_5 gnd vdd FILL
XFILL_34_DFFSR_198 gnd vdd FILL
XFILL_11_AOI21X1_65 gnd vdd FILL
XFILL_38_DFFSR_120 gnd vdd FILL
XFILL_11_AOI21X1_76 gnd vdd FILL
XFILL_38_DFFSR_131 gnd vdd FILL
XFILL_38_DFFSR_142 gnd vdd FILL
XFILL_38_DFFSR_153 gnd vdd FILL
XFILL_58_DFFSR_3 gnd vdd FILL
XFILL_38_DFFSR_164 gnd vdd FILL
XFILL_30_NOR3X1_11 gnd vdd FILL
XFILL_38_DFFSR_175 gnd vdd FILL
XFILL_2_INVX1_19 gnd vdd FILL
XFILL_38_DFFSR_186 gnd vdd FILL
XFILL_30_NOR3X1_22 gnd vdd FILL
XFILL_38_DFFSR_197 gnd vdd FILL
XFILL_30_NOR3X1_33 gnd vdd FILL
XFILL_80_DFFSR_200 gnd vdd FILL
XFILL_30_NOR3X1_44 gnd vdd FILL
XFILL_80_DFFSR_211 gnd vdd FILL
XFILL_80_DFFSR_222 gnd vdd FILL
XFILL_2_1 gnd vdd FILL
XFILL_80_DFFSR_233 gnd vdd FILL
XFILL_80_DFFSR_244 gnd vdd FILL
XFILL_80_DFFSR_255 gnd vdd FILL
XFILL_80_DFFSR_266 gnd vdd FILL
XFILL_84_DFFSR_210 gnd vdd FILL
XFILL_84_DFFSR_221 gnd vdd FILL
XFILL_11_AOI21X1_6 gnd vdd FILL
XFILL_0_BUFX4_17 gnd vdd FILL
XFILL_37_6_2 gnd vdd FILL
XFILL_84_DFFSR_232 gnd vdd FILL
XFILL_84_DFFSR_243 gnd vdd FILL
XFILL_42_DFFSR_9 gnd vdd FILL
XFILL_0_BUFX4_28 gnd vdd FILL
XFILL_84_DFFSR_254 gnd vdd FILL
XFILL_0_BUFX4_39 gnd vdd FILL
XFILL_44_1 gnd vdd FILL
XFILL_36_1_1 gnd vdd FILL
XFILL_84_DFFSR_265 gnd vdd FILL
XFILL_6_CLKBUF1_30 gnd vdd FILL
XFILL_6_CLKBUF1_41 gnd vdd FILL
XFILL_14_MUX2X1_104 gnd vdd FILL
XFILL_14_MUX2X1_115 gnd vdd FILL
XFILL_15_AOI21X1_5 gnd vdd FILL
XFILL_14_MUX2X1_126 gnd vdd FILL
XFILL_0_INVX1_160 gnd vdd FILL
XFILL_14_MUX2X1_137 gnd vdd FILL
XFILL_14_MUX2X1_148 gnd vdd FILL
XFILL_0_INVX1_171 gnd vdd FILL
XFILL_0_INVX1_182 gnd vdd FILL
XFILL_14_MUX2X1_159 gnd vdd FILL
XFILL_1_AOI21X1_60 gnd vdd FILL
XFILL_0_INVX1_193 gnd vdd FILL
XFILL_1_AOI21X1_71 gnd vdd FILL
XFILL_11_OAI22X1_40 gnd vdd FILL
XFILL_11_OAI22X1_51 gnd vdd FILL
XFILL_15_OAI21X1_20 gnd vdd FILL
XFILL_15_OAI21X1_31 gnd vdd FILL
XFILL_4_INVX1_170 gnd vdd FILL
XFILL_15_OAI21X1_42 gnd vdd FILL
XFILL_20_5_2 gnd vdd FILL
XFILL_4_INVX1_181 gnd vdd FILL
XFILL_4_INVX1_192 gnd vdd FILL
XFILL_4_NOR2X1_170 gnd vdd FILL
XFILL_4_NOR2X1_181 gnd vdd FILL
XFILL_4_NOR2X1_192 gnd vdd FILL
XFILL_26_DFFSR_19 gnd vdd FILL
XFILL_66_DFFSR_18 gnd vdd FILL
XFILL_66_DFFSR_29 gnd vdd FILL
XFILL_21_MUX2X1_150 gnd vdd FILL
XFILL_21_MUX2X1_161 gnd vdd FILL
XFILL_4_MUX2X1_110 gnd vdd FILL
XFILL_21_MUX2X1_172 gnd vdd FILL
XFILL_4_MUX2X1_121 gnd vdd FILL
XNAND3X1_17 NAND3X1_17/A INVX1_129/Y NAND3X1_17/C gnd NOR3X1_44/C vdd NAND3X1
XFILL_21_MUX2X1_183 gnd vdd FILL
XFILL_21_MUX2X1_194 gnd vdd FILL
XNAND3X1_28 OAI21X1_48/A OAI21X1_41/A AND2X2_7/Y gnd NAND3X1_29/C vdd NAND3X1
XFILL_4_MUX2X1_132 gnd vdd FILL
XNAND3X1_39 DFFSR_1/D NAND3X1_39/B OAI21X1_45/Y gnd NOR3X1_9/C vdd NAND3X1
XFILL_4_MUX2X1_143 gnd vdd FILL
XFILL_4_MUX2X1_154 gnd vdd FILL
XFILL_4_MUX2X1_165 gnd vdd FILL
XFILL_4_BUFX4_8 gnd vdd FILL
XFILL_4_MUX2X1_176 gnd vdd FILL
XFILL_7_NAND3X1_109 gnd vdd FILL
XFILL_35_DFFSR_17 gnd vdd FILL
XFILL_4_MUX2X1_187 gnd vdd FILL
XFILL_35_DFFSR_28 gnd vdd FILL
XNOR2X1_17 NOR2X1_7/B INVX1_8/Y gnd NOR2X1_19/B vdd NOR2X1
XFILL_35_DFFSR_39 gnd vdd FILL
XNOR2X1_28 NOR2X1_28/A NOR2X1_28/B gnd NOR2X1_28/Y vdd NOR2X1
XFILL_28_6_2 gnd vdd FILL
XFILL_3_6_2 gnd vdd FILL
XFILL_51_DFFSR_210 gnd vdd FILL
XNOR2X1_39 NOR2X1_39/A NOR2X1_39/B gnd NOR2X1_39/Y vdd NOR2X1
XFILL_51_DFFSR_221 gnd vdd FILL
XFILL_27_1_1 gnd vdd FILL
XFILL_2_1_1 gnd vdd FILL
XFILL_51_DFFSR_232 gnd vdd FILL
XFILL_51_DFFSR_243 gnd vdd FILL
XFILL_51_DFFSR_254 gnd vdd FILL
XFILL_75_DFFSR_16 gnd vdd FILL
XFILL_75_DFFSR_27 gnd vdd FILL
XFILL_51_DFFSR_265 gnd vdd FILL
XFILL_75_DFFSR_38 gnd vdd FILL
XFILL_75_DFFSR_49 gnd vdd FILL
XFILL_18_MUX2X1_6 gnd vdd FILL
XFILL_55_DFFSR_220 gnd vdd FILL
XFILL_11_NAND3X1_100 gnd vdd FILL
XFILL_55_DFFSR_231 gnd vdd FILL
XFILL_55_DFFSR_242 gnd vdd FILL
XFILL_11_NAND3X1_111 gnd vdd FILL
XFILL_55_DFFSR_253 gnd vdd FILL
XFILL_11_NAND3X1_122 gnd vdd FILL
XFILL_55_DFFSR_264 gnd vdd FILL
XFILL_55_DFFSR_275 gnd vdd FILL
XFILL_10_CLKBUF1_5 gnd vdd FILL
XFILL_9_BUFX4_50 gnd vdd FILL
XFILL_9_BUFX4_61 gnd vdd FILL
XFILL_11_5_2 gnd vdd FILL
XFILL_44_DFFSR_15 gnd vdd FILL
XFILL_0_BUFX2_4 gnd vdd FILL
XFILL_82_DFFSR_120 gnd vdd FILL
XFILL_44_DFFSR_26 gnd vdd FILL
XFILL_9_BUFX4_72 gnd vdd FILL
XFILL_82_DFFSR_131 gnd vdd FILL
XFILL_9_BUFX4_83 gnd vdd FILL
XFILL_44_DFFSR_37 gnd vdd FILL
XFILL_59_DFFSR_230 gnd vdd FILL
XFILL_10_0_1 gnd vdd FILL
XFILL_82_DFFSR_142 gnd vdd FILL
XFILL_44_DFFSR_48 gnd vdd FILL
XFILL_9_BUFX4_94 gnd vdd FILL
XFILL_82_DFFSR_153 gnd vdd FILL
XFILL_59_DFFSR_241 gnd vdd FILL
XFILL_59_DFFSR_252 gnd vdd FILL
XFILL_44_DFFSR_59 gnd vdd FILL
XFILL_59_DFFSR_263 gnd vdd FILL
XFILL_82_DFFSR_164 gnd vdd FILL
XFILL_59_DFFSR_274 gnd vdd FILL
XFILL_82_DFFSR_175 gnd vdd FILL
XFILL_14_CLKBUF1_4 gnd vdd FILL
XFILL_2_DFFSR_201 gnd vdd FILL
XFILL_82_DFFSR_186 gnd vdd FILL
XFILL_82_DFFSR_197 gnd vdd FILL
XFILL_2_DFFSR_212 gnd vdd FILL
XFILL_84_DFFSR_14 gnd vdd FILL
XFILL_2_DFFSR_223 gnd vdd FILL
XFILL_84_DFFSR_25 gnd vdd FILL
XFILL_7_NAND3X1_13 gnd vdd FILL
XFILL_86_DFFSR_130 gnd vdd FILL
XFILL_2_DFFSR_234 gnd vdd FILL
XFILL_84_DFFSR_36 gnd vdd FILL
XFILL_7_NAND3X1_24 gnd vdd FILL
XFILL_2_DFFSR_245 gnd vdd FILL
XFILL_7_NAND3X1_35 gnd vdd FILL
XFILL_86_DFFSR_141 gnd vdd FILL
XFILL_2_NAND3X1_105 gnd vdd FILL
XFILL_84_DFFSR_47 gnd vdd FILL
XFILL_86_DFFSR_152 gnd vdd FILL
XFILL_84_DFFSR_58 gnd vdd FILL
XFILL_2_DFFSR_256 gnd vdd FILL
XFILL_7_NAND3X1_46 gnd vdd FILL
XFILL_2_DFFSR_267 gnd vdd FILL
XFILL_2_NAND3X1_116 gnd vdd FILL
XFILL_13_DFFSR_14 gnd vdd FILL
XFILL_86_DFFSR_163 gnd vdd FILL
XFILL_7_NAND3X1_57 gnd vdd FILL
XFILL_84_DFFSR_69 gnd vdd FILL
XFILL_13_DFFSR_25 gnd vdd FILL
XFILL_2_NAND3X1_127 gnd vdd FILL
XFILL_86_DFFSR_174 gnd vdd FILL
XFILL_18_CLKBUF1_3 gnd vdd FILL
XFILL_7_NAND3X1_68 gnd vdd FILL
XFILL_13_DFFSR_36 gnd vdd FILL
XFILL_6_DFFSR_200 gnd vdd FILL
XFILL_7_NAND3X1_79 gnd vdd FILL
XFILL_86_DFFSR_185 gnd vdd FILL
XFILL_13_DFFSR_47 gnd vdd FILL
XFILL_6_DFFSR_211 gnd vdd FILL
XFILL_13_DFFSR_58 gnd vdd FILL
XFILL_86_DFFSR_196 gnd vdd FILL
XFILL_6_DFFSR_222 gnd vdd FILL
XFILL_37_DFFSR_209 gnd vdd FILL
XFILL_13_DFFSR_69 gnd vdd FILL
XFILL_6_DFFSR_233 gnd vdd FILL
XFILL_6_DFFSR_244 gnd vdd FILL
XFILL_53_DFFSR_13 gnd vdd FILL
XFILL_6_DFFSR_255 gnd vdd FILL
XFILL_6_DFFSR_266 gnd vdd FILL
XFILL_53_DFFSR_24 gnd vdd FILL
XFILL_53_DFFSR_35 gnd vdd FILL
XFILL_53_DFFSR_46 gnd vdd FILL
XFILL_53_DFFSR_57 gnd vdd FILL
XFILL_64_DFFSR_109 gnd vdd FILL
XFILL_53_DFFSR_68 gnd vdd FILL
XFILL_53_DFFSR_79 gnd vdd FILL
XMUX2X1_13 MUX2X1_4/B INVX1_46/Y NOR2X1_2/B gnd MUX2X1_13/Y vdd MUX2X1
XFILL_19_6_2 gnd vdd FILL
XFILL_0_NAND2X1_15 gnd vdd FILL
XFILL_0_NAND2X1_26 gnd vdd FILL
XMUX2X1_24 BUFX4_66/Y INVX1_79/Y NOR2X1_2/B gnd MUX2X1_24/Y vdd MUX2X1
XFILL_24_DFFSR_6 gnd vdd FILL
XMUX2X1_35 BUFX4_93/Y INVX1_90/Y NOR2X1_2/B gnd MUX2X1_35/Y vdd MUX2X1
XFILL_18_1_1 gnd vdd FILL
XFILL_0_NAND2X1_37 gnd vdd FILL
XFILL_68_DFFSR_108 gnd vdd FILL
XFILL_22_DFFSR_12 gnd vdd FILL
XFILL_0_NAND2X1_48 gnd vdd FILL
XNOR2X1_107 OAI21X1_32/Y OAI21X1_31/Y gnd NOR2X1_107/Y vdd NOR2X1
XMUX2X1_46 MUX2X1_4/B NOR3X1_45/A NOR2X1_46/B gnd MUX2X1_46/Y vdd MUX2X1
XNOR2X1_118 INVX2_4/Y OAI21X1_48/A gnd OAI21X1_45/B vdd NOR2X1
XFILL_0_NAND2X1_59 gnd vdd FILL
XMUX2X1_57 MUX2X1_9/A NOR3X1_15/A NOR2X1_46/B gnd MUX2X1_57/Y vdd MUX2X1
XFILL_22_DFFSR_23 gnd vdd FILL
XNOR2X1_129 NOR2X1_27/A INVX4_1/Y gnd AOI21X1_7/B vdd NOR2X1
XMUX2X1_68 BUFX4_93/Y NOR3X1_40/A NOR2X1_46/B gnd MUX2X1_68/Y vdd MUX2X1
XFILL_68_DFFSR_119 gnd vdd FILL
XFILL_81_DFFSR_7 gnd vdd FILL
XMUX2X1_79 BUFX4_81/Y OAI21X1_4/A NOR2X1_57/Y gnd MUX2X1_79/Y vdd MUX2X1
XFILL_22_DFFSR_34 gnd vdd FILL
XFILL_22_DFFSR_45 gnd vdd FILL
XFILL_22_DFFSR_56 gnd vdd FILL
XFILL_11_OAI21X1_9 gnd vdd FILL
XFILL_61_4_2 gnd vdd FILL
XFILL_22_DFFSR_67 gnd vdd FILL
XFILL_0_INVX2_4 gnd vdd FILL
XFILL_22_DFFSR_78 gnd vdd FILL
XFILL_22_DFFSR_89 gnd vdd FILL
XFILL_23_6 gnd vdd FILL
XFILL_62_DFFSR_11 gnd vdd FILL
XFILL_10_MUX2X1_190 gnd vdd FILL
XFILL_62_DFFSR_22 gnd vdd FILL
XFILL_62_DFFSR_33 gnd vdd FILL
XFILL_22_DFFSR_220 gnd vdd FILL
XFILL_3_AOI22X1_5 gnd vdd FILL
XFILL_16_5 gnd vdd FILL
XFILL_62_DFFSR_44 gnd vdd FILL
XFILL_62_DFFSR_55 gnd vdd FILL
XFILL_15_OAI21X1_8 gnd vdd FILL
XFILL_22_DFFSR_231 gnd vdd FILL
XFILL_22_DFFSR_242 gnd vdd FILL
XFILL_62_DFFSR_66 gnd vdd FILL
XFILL_62_DFFSR_77 gnd vdd FILL
XFILL_22_DFFSR_253 gnd vdd FILL
XFILL_62_DFFSR_88 gnd vdd FILL
XFILL_22_DFFSR_264 gnd vdd FILL
XFILL_22_DFFSR_275 gnd vdd FILL
XFILL_62_DFFSR_99 gnd vdd FILL
XFILL_3_INVX1_204 gnd vdd FILL
XFILL_3_INVX1_215 gnd vdd FILL
XFILL_26_CLKBUF1_14 gnd vdd FILL
XFILL_5_DFFSR_13 gnd vdd FILL
XDFFSR_5 DFFSR_5/Q DFFSR_5/CLK DFFSR_5/R vdd DFFSR_5/D gnd vdd DFFSR
XFILL_26_CLKBUF1_25 gnd vdd FILL
XFILL_5_DFFSR_24 gnd vdd FILL
XFILL_3_INVX1_226 gnd vdd FILL
XFILL_26_CLKBUF1_36 gnd vdd FILL
XFILL_26_DFFSR_230 gnd vdd FILL
XFILL_7_AOI22X1_4 gnd vdd FILL
XFILL_5_DFFSR_35 gnd vdd FILL
XFILL_31_DFFSR_10 gnd vdd FILL
XFILL_31_DFFSR_21 gnd vdd FILL
XFILL_5_DFFSR_46 gnd vdd FILL
XFILL_26_DFFSR_241 gnd vdd FILL
XFILL_5_DFFSR_57 gnd vdd FILL
XFILL_26_DFFSR_252 gnd vdd FILL
XFILL_31_DFFSR_32 gnd vdd FILL
XFILL_31_DFFSR_43 gnd vdd FILL
XFILL_5_DFFSR_68 gnd vdd FILL
XFILL_26_DFFSR_263 gnd vdd FILL
XFILL_26_DFFSR_274 gnd vdd FILL
XFILL_9_CLKBUF1_18 gnd vdd FILL
XFILL_5_DFFSR_79 gnd vdd FILL
XFILL_9_CLKBUF1_29 gnd vdd FILL
XFILL_7_INVX1_203 gnd vdd FILL
XFILL_31_DFFSR_54 gnd vdd FILL
XFILL_23_MUX2X1_19 gnd vdd FILL
XFILL_31_DFFSR_65 gnd vdd FILL
XFILL_7_INVX1_214 gnd vdd FILL
XFILL_31_DFFSR_76 gnd vdd FILL
XFILL_7_INVX1_225 gnd vdd FILL
XFILL_4_AOI21X1_15 gnd vdd FILL
XFILL_31_DFFSR_87 gnd vdd FILL
XFILL_53_DFFSR_130 gnd vdd FILL
XFILL_31_DFFSR_98 gnd vdd FILL
XFILL_4_AOI21X1_26 gnd vdd FILL
XFILL_53_DFFSR_141 gnd vdd FILL
XFILL_53_DFFSR_152 gnd vdd FILL
XFILL_71_DFFSR_20 gnd vdd FILL
XFILL_4_AOI21X1_37 gnd vdd FILL
XFILL_71_DFFSR_31 gnd vdd FILL
XFILL_4_AOI21X1_48 gnd vdd FILL
XFILL_4_AOI21X1_59 gnd vdd FILL
XFILL_71_DFFSR_42 gnd vdd FILL
XFILL_53_DFFSR_163 gnd vdd FILL
XFILL_53_DFFSR_174 gnd vdd FILL
XFILL_14_OAI22X1_17 gnd vdd FILL
XFILL_71_DFFSR_53 gnd vdd FILL
XFILL_14_OAI22X1_28 gnd vdd FILL
XFILL_53_DFFSR_185 gnd vdd FILL
XFILL_71_DFFSR_64 gnd vdd FILL
XFILL_14_OAI22X1_39 gnd vdd FILL
XFILL_53_DFFSR_196 gnd vdd FILL
XFILL_7_NOR2X1_103 gnd vdd FILL
XFILL_71_DFFSR_75 gnd vdd FILL
XFILL_71_DFFSR_86 gnd vdd FILL
XFILL_7_NOR2X1_114 gnd vdd FILL
XFILL_71_DFFSR_97 gnd vdd FILL
XFILL_7_NOR2X1_125 gnd vdd FILL
XFILL_57_DFFSR_140 gnd vdd FILL
XFILL_57_DFFSR_151 gnd vdd FILL
XFILL_7_NOR2X1_136 gnd vdd FILL
XFILL_57_DFFSR_162 gnd vdd FILL
XFILL_7_NOR2X1_147 gnd vdd FILL
XFILL_7_NOR2X1_158 gnd vdd FILL
XFILL_0_DFFSR_100 gnd vdd FILL
XFILL_57_DFFSR_173 gnd vdd FILL
XFILL_7_NOR2X1_169 gnd vdd FILL
XFILL_57_DFFSR_184 gnd vdd FILL
XNAND2X1_50 BUFX4_89/Y AND2X2_1/Y gnd OAI21X1_2/B vdd NAND2X1
XFILL_13_NAND3X1_60 gnd vdd FILL
XFILL_57_DFFSR_195 gnd vdd FILL
XFILL_0_DFFSR_111 gnd vdd FILL
XNAND2X1_61 NOR2X1_63/Y NOR2X1_64/Y gnd NOR3X1_18/B vdd NAND2X1
XFILL_31_DFFSR_109 gnd vdd FILL
XFILL_13_NAND3X1_71 gnd vdd FILL
XNAND2X1_72 INVX1_65/A NOR2X1_69/Y gnd NAND2X1_72/Y vdd NAND2X1
XFILL_40_DFFSR_30 gnd vdd FILL
XFILL_0_DFFSR_122 gnd vdd FILL
XFILL_0_DFFSR_133 gnd vdd FILL
XFILL_13_NAND3X1_82 gnd vdd FILL
XFILL_40_DFFSR_41 gnd vdd FILL
XFILL_11_NOR3X1_5 gnd vdd FILL
XFILL_0_DFFSR_144 gnd vdd FILL
XNAND2X1_83 INVX2_3/A BUFX2_7/A gnd OAI21X1_46/B vdd NAND2X1
XFILL_40_DFFSR_52 gnd vdd FILL
XFILL_40_DFFSR_63 gnd vdd FILL
XFILL_13_NAND3X1_93 gnd vdd FILL
XFILL_0_DFFSR_155 gnd vdd FILL
XNAND2X1_94 NAND3X1_43/B OAI21X1_42/Y gnd DFFSR_112/D vdd NAND2X1
XFILL_40_DFFSR_74 gnd vdd FILL
XFILL_0_DFFSR_166 gnd vdd FILL
XFILL_0_DFFSR_177 gnd vdd FILL
XFILL_40_DFFSR_85 gnd vdd FILL
XFILL_40_DFFSR_96 gnd vdd FILL
XFILL_0_DFFSR_188 gnd vdd FILL
XFILL_4_DFFSR_110 gnd vdd FILL
XFILL_0_DFFSR_199 gnd vdd FILL
XFILL_35_DFFSR_108 gnd vdd FILL
XFILL_52_4_2 gnd vdd FILL
XFILL_4_DFFSR_121 gnd vdd FILL
XFILL_80_DFFSR_40 gnd vdd FILL
XFILL_4_DFFSR_132 gnd vdd FILL
XFILL_35_DFFSR_119 gnd vdd FILL
XFILL_80_DFFSR_51 gnd vdd FILL
XFILL_4_DFFSR_143 gnd vdd FILL
XFILL_4_DFFSR_154 gnd vdd FILL
XFILL_80_DFFSR_62 gnd vdd FILL
XFILL_80_DFFSR_73 gnd vdd FILL
XFILL_4_DFFSR_165 gnd vdd FILL
XFILL_80_DFFSR_84 gnd vdd FILL
XFILL_4_DFFSR_176 gnd vdd FILL
XFILL_80_DFFSR_95 gnd vdd FILL
XFILL_4_DFFSR_187 gnd vdd FILL
XFILL_4_DFFSR_198 gnd vdd FILL
XFILL_39_DFFSR_107 gnd vdd FILL
XFILL_7_MUX2X1_109 gnd vdd FILL
XFILL_8_DFFSR_120 gnd vdd FILL
XFILL_8_DFFSR_131 gnd vdd FILL
XFILL_39_DFFSR_118 gnd vdd FILL
XFILL_8_DFFSR_142 gnd vdd FILL
XFILL_12_MUX2X1_40 gnd vdd FILL
XFILL_39_DFFSR_129 gnd vdd FILL
XFILL_8_DFFSR_153 gnd vdd FILL
XFILL_12_MUX2X1_51 gnd vdd FILL
XFILL_8_BUFX4_9 gnd vdd FILL
XFILL_12_MUX2X1_62 gnd vdd FILL
XFILL_4_OAI22X1_12 gnd vdd FILL
XFILL_8_DFFSR_164 gnd vdd FILL
XFILL_20_NOR3X1_3 gnd vdd FILL
XFILL_4_OAI22X1_23 gnd vdd FILL
XFILL_12_MUX2X1_73 gnd vdd FILL
XFILL_0_NOR3X1_11 gnd vdd FILL
XFILL_8_DFFSR_175 gnd vdd FILL
XFILL_12_MUX2X1_84 gnd vdd FILL
XFILL_8_DFFSR_186 gnd vdd FILL
XFILL_4_OAI22X1_34 gnd vdd FILL
XFILL_0_NOR3X1_22 gnd vdd FILL
XFILL_8_DFFSR_197 gnd vdd FILL
XFILL_0_NOR3X1_33 gnd vdd FILL
XFILL_12_MUX2X1_95 gnd vdd FILL
XFILL_4_OAI22X1_45 gnd vdd FILL
XFILL_8_OAI21X1_14 gnd vdd FILL
XFILL_0_NOR3X1_44 gnd vdd FILL
XFILL_8_OAI21X1_25 gnd vdd FILL
XFILL_8_OAI21X1_36 gnd vdd FILL
XFILL_81_DFFSR_209 gnd vdd FILL
XFILL_8_OAI21X1_47 gnd vdd FILL
XFILL_16_MUX2X1_50 gnd vdd FILL
XFILL_16_MUX2X1_61 gnd vdd FILL
XFILL_16_MUX2X1_72 gnd vdd FILL
XFILL_4_NOR3X1_10 gnd vdd FILL
XFILL_16_MUX2X1_83 gnd vdd FILL
XFILL_4_NOR3X1_21 gnd vdd FILL
XFILL_16_MUX2X1_94 gnd vdd FILL
XFILL_4_NOR3X1_32 gnd vdd FILL
XFILL_4_NOR3X1_43 gnd vdd FILL
XFILL_85_DFFSR_208 gnd vdd FILL
XFILL_1_NOR2X1_203 gnd vdd FILL
XFILL_20_DFFSR_130 gnd vdd FILL
XFILL_85_DFFSR_219 gnd vdd FILL
XFILL_20_DFFSR_141 gnd vdd FILL
XFILL_20_DFFSR_152 gnd vdd FILL
XFILL_7_NAND2X1_90 gnd vdd FILL
XFILL_20_DFFSR_163 gnd vdd FILL
XFILL_3_NOR3X1_4 gnd vdd FILL
XFILL_8_NOR3X1_20 gnd vdd FILL
XFILL_20_DFFSR_174 gnd vdd FILL
XFILL_8_NOR3X1_31 gnd vdd FILL
XFILL_1_INVX1_103 gnd vdd FILL
XFILL_59_0_1 gnd vdd FILL
XFILL_8_NOR3X1_42 gnd vdd FILL
XFILL_20_DFFSR_185 gnd vdd FILL
XFILL_1_INVX1_114 gnd vdd FILL
XFILL_15_CLKBUF1_10 gnd vdd FILL
XFILL_20_DFFSR_196 gnd vdd FILL
XFILL_1_INVX1_125 gnd vdd FILL
XFILL_15_CLKBUF1_21 gnd vdd FILL
XFILL_4_BUFX2_5 gnd vdd FILL
XFILL_1_INVX1_136 gnd vdd FILL
XFILL_15_CLKBUF1_32 gnd vdd FILL
XFILL_1_INVX1_147 gnd vdd FILL
XFILL_24_DFFSR_140 gnd vdd FILL
XFILL_24_DFFSR_151 gnd vdd FILL
XFILL_1_INVX1_158 gnd vdd FILL
XFILL_24_DFFSR_162 gnd vdd FILL
XFILL_1_INVX1_169 gnd vdd FILL
XFILL_5_INVX1_102 gnd vdd FILL
XFILL_10_AOI21X1_40 gnd vdd FILL
XFILL_24_DFFSR_173 gnd vdd FILL
XFILL_24_DFFSR_184 gnd vdd FILL
XFILL_10_AOI21X1_51 gnd vdd FILL
XFILL_5_INVX1_113 gnd vdd FILL
XFILL_10_AOI21X1_62 gnd vdd FILL
XFILL_24_DFFSR_195 gnd vdd FILL
XFILL_5_INVX1_124 gnd vdd FILL
XFILL_10_AOI21X1_73 gnd vdd FILL
XFILL_5_INVX1_135 gnd vdd FILL
XFILL_5_INVX1_146 gnd vdd FILL
XFILL_5_INVX1_157 gnd vdd FILL
XFILL_1_DFFSR_50 gnd vdd FILL
XFILL_63_DFFSR_4 gnd vdd FILL
XFILL_28_DFFSR_150 gnd vdd FILL
XFILL_1_DFFSR_61 gnd vdd FILL
XFILL_28_DFFSR_161 gnd vdd FILL
XFILL_5_INVX1_168 gnd vdd FILL
XFILL_1_DFFSR_72 gnd vdd FILL
XFILL_1_DFFSR_83 gnd vdd FILL
XFILL_43_4_2 gnd vdd FILL
XFILL_28_DFFSR_172 gnd vdd FILL
XFILL_5_INVX1_179 gnd vdd FILL
XFILL_1_DFFSR_94 gnd vdd FILL
XFILL_2_OR2X2_1 gnd vdd FILL
XFILL_28_DFFSR_183 gnd vdd FILL
XFILL_28_DFFSR_194 gnd vdd FILL
XFILL_20_NOR3X1_30 gnd vdd FILL
XFILL_20_NOR3X1_41 gnd vdd FILL
XFILL_20_NOR3X1_52 gnd vdd FILL
XFILL_12_NAND3X1_101 gnd vdd FILL
XFILL_70_DFFSR_230 gnd vdd FILL
XFILL_70_DFFSR_241 gnd vdd FILL
XFILL_12_NAND3X1_112 gnd vdd FILL
XFILL_12_NAND3X1_123 gnd vdd FILL
XFILL_70_DFFSR_252 gnd vdd FILL
XFILL_70_DFFSR_263 gnd vdd FILL
XFILL_70_DFFSR_274 gnd vdd FILL
XFILL_24_NOR3X1_40 gnd vdd FILL
XFILL_24_NOR3X1_51 gnd vdd FILL
XFILL_3_OAI22X1_8 gnd vdd FILL
XFILL_74_DFFSR_240 gnd vdd FILL
XFILL_74_DFFSR_251 gnd vdd FILL
XFILL_74_DFFSR_262 gnd vdd FILL
XFILL_74_DFFSR_273 gnd vdd FILL
XFILL_28_DFFSR_7 gnd vdd FILL
XFILL_28_NOR3X1_50 gnd vdd FILL
XFILL_85_DFFSR_8 gnd vdd FILL
XFILL_13_MUX2X1_101 gnd vdd FILL
XFILL_13_MUX2X1_112 gnd vdd FILL
XFILL_13_MUX2X1_123 gnd vdd FILL
XFILL_7_OAI22X1_7 gnd vdd FILL
XFILL_4_INVX2_5 gnd vdd FILL
XFILL_13_MUX2X1_134 gnd vdd FILL
XFILL_3_NAND3X1_106 gnd vdd FILL
XFILL_13_MUX2X1_145 gnd vdd FILL
XFILL_3_NAND3X1_117 gnd vdd FILL
XFILL_13_MUX2X1_156 gnd vdd FILL
XFILL_78_DFFSR_250 gnd vdd FILL
XFILL_3_NAND3X1_128 gnd vdd FILL
XFILL_13_MUX2X1_167 gnd vdd FILL
XFILL_78_DFFSR_261 gnd vdd FILL
XFILL_78_DFFSR_272 gnd vdd FILL
XFILL_33_CLKBUF1_2 gnd vdd FILL
XFILL_13_MUX2X1_178 gnd vdd FILL
XFILL_13_MUX2X1_189 gnd vdd FILL
XFILL_52_DFFSR_208 gnd vdd FILL
XFILL_52_DFFSR_219 gnd vdd FILL
XFILL_14_OAI21X1_50 gnd vdd FILL
XFILL_2_INVX1_3 gnd vdd FILL
XFILL_56_DFFSR_207 gnd vdd FILL
XFILL_56_DFFSR_218 gnd vdd FILL
XFILL_56_DFFSR_229 gnd vdd FILL
XFILL_62_7_0 gnd vdd FILL
XFILL_83_DFFSR_107 gnd vdd FILL
XFILL_34_4_2 gnd vdd FILL
XFILL_83_DFFSR_118 gnd vdd FILL
XFILL_83_DFFSR_129 gnd vdd FILL
XFILL_21_3 gnd vdd FILL
XFILL_87_DFFSR_106 gnd vdd FILL
XFILL_20_MUX2X1_180 gnd vdd FILL
XFILL_87_DFFSR_117 gnd vdd FILL
XFILL_14_2 gnd vdd FILL
XFILL_20_MUX2X1_191 gnd vdd FILL
XFILL_14_BUFX4_11 gnd vdd FILL
XFILL_3_MUX2X1_140 gnd vdd FILL
XFILL_87_DFFSR_128 gnd vdd FILL
XFILL_14_BUFX4_22 gnd vdd FILL
XFILL_87_DFFSR_139 gnd vdd FILL
XFILL_3_MUX2X1_151 gnd vdd FILL
XFILL_3_MUX2X1_162 gnd vdd FILL
XFILL_14_BUFX4_33 gnd vdd FILL
XFILL_3_MUX2X1_173 gnd vdd FILL
XFILL_14_BUFX4_44 gnd vdd FILL
XFILL_3_MUX2X1_184 gnd vdd FILL
XDFFSR_201 INVX1_93/A DFFSR_45/CLK BUFX4_13/Y vdd MUX2X1_80/Y gnd vdd DFFSR
XFILL_14_BUFX4_55 gnd vdd FILL
XDFFSR_212 INVX1_87/A DFFSR_79/CLK DFFSR_79/R vdd MUX2X1_74/Y gnd vdd DFFSR
XFILL_14_BUFX4_66 gnd vdd FILL
XDFFSR_223 INVX1_72/A CLKBUF1_26/Y DFFSR_25/R vdd MUX2X1_59/Y gnd vdd DFFSR
XFILL_14_BUFX4_77 gnd vdd FILL
XFILL_7_DFFSR_209 gnd vdd FILL
XDFFSR_234 INVX1_65/A DFFSR_4/CLK DFFSR_23/R vdd MUX2X1_52/Y gnd vdd DFFSR
XFILL_4_NAND3X1_9 gnd vdd FILL
XFILL_14_BUFX4_88 gnd vdd FILL
XFILL_14_BUFX4_99 gnd vdd FILL
XDFFSR_245 INVX1_50/A DFFSR_39/CLK DFFSR_45/R vdd MUX2X1_37/Y gnd vdd DFFSR
XDFFSR_256 INVX1_44/A DFFSR_8/CLK DFFSR_8/R vdd MUX2X1_31/Y gnd vdd DFFSR
XDFFSR_267 NOR2X1_8/A DFFSR_1/CLK BUFX4_54/Y vdd DFFSR_267/D gnd vdd DFFSR
XFILL_41_DFFSR_240 gnd vdd FILL
XFILL_41_DFFSR_251 gnd vdd FILL
XFILL_41_DFFSR_262 gnd vdd FILL
XFILL_41_DFFSR_273 gnd vdd FILL
XFILL_8_NAND3X1_8 gnd vdd FILL
XFILL_45_DFFSR_250 gnd vdd FILL
XFILL_45_DFFSR_261 gnd vdd FILL
XFILL_45_DFFSR_272 gnd vdd FILL
XFILL_9_AND2X2_4 gnd vdd FILL
XFILL_72_DFFSR_150 gnd vdd FILL
XFILL_72_DFFSR_161 gnd vdd FILL
XFILL_49_DFFSR_260 gnd vdd FILL
XFILL_49_DFFSR_271 gnd vdd FILL
XFILL_72_DFFSR_172 gnd vdd FILL
XFILL_72_DFFSR_183 gnd vdd FILL
XFILL_72_DFFSR_194 gnd vdd FILL
XFILL_23_DFFSR_207 gnd vdd FILL
XFILL_23_DFFSR_218 gnd vdd FILL
XFILL_6_NAND3X1_10 gnd vdd FILL
XFILL_6_NAND3X1_21 gnd vdd FILL
XFILL_6_NAND3X1_32 gnd vdd FILL
XFILL_23_DFFSR_229 gnd vdd FILL
XFILL_53_7_0 gnd vdd FILL
XFILL_6_NAND3X1_43 gnd vdd FILL
XFILL_76_DFFSR_160 gnd vdd FILL
XFILL_25_4_2 gnd vdd FILL
XFILL_6_NAND3X1_54 gnd vdd FILL
XFILL_0_4_2 gnd vdd FILL
XFILL_45_DFFSR_1 gnd vdd FILL
XFILL_76_DFFSR_171 gnd vdd FILL
XFILL_6_BUFX4_10 gnd vdd FILL
XFILL_6_NAND3X1_65 gnd vdd FILL
XFILL_6_NAND3X1_76 gnd vdd FILL
XFILL_76_DFFSR_182 gnd vdd FILL
XFILL_6_NAND3X1_87 gnd vdd FILL
XFILL_76_DFFSR_193 gnd vdd FILL
XFILL_6_BUFX4_21 gnd vdd FILL
XFILL_27_DFFSR_206 gnd vdd FILL
XFILL_50_DFFSR_107 gnd vdd FILL
XFILL_6_BUFX4_32 gnd vdd FILL
XFILL_6_NAND3X1_98 gnd vdd FILL
XFILL_27_DFFSR_217 gnd vdd FILL
XFILL_6_BUFX4_43 gnd vdd FILL
XFILL_50_DFFSR_118 gnd vdd FILL
XFILL_6_BUFX4_54 gnd vdd FILL
XFILL_27_DFFSR_228 gnd vdd FILL
XFILL_50_DFFSR_129 gnd vdd FILL
XFILL_6_BUFX4_65 gnd vdd FILL
XFILL_41_DFFSR_19 gnd vdd FILL
XFILL_27_DFFSR_239 gnd vdd FILL
XFILL_6_BUFX4_76 gnd vdd FILL
XFILL_6_BUFX4_87 gnd vdd FILL
XFILL_6_BUFX4_98 gnd vdd FILL
XFILL_54_DFFSR_106 gnd vdd FILL
XFILL_8_BUFX2_6 gnd vdd FILL
XFILL_54_DFFSR_117 gnd vdd FILL
XFILL_54_DFFSR_128 gnd vdd FILL
XFILL_54_DFFSR_139 gnd vdd FILL
XFILL_81_DFFSR_18 gnd vdd FILL
XFILL_13_AOI21X1_17 gnd vdd FILL
XFILL_81_DFFSR_29 gnd vdd FILL
XFILL_13_AOI21X1_28 gnd vdd FILL
XFILL_13_AOI21X1_39 gnd vdd FILL
XFILL_58_DFFSR_105 gnd vdd FILL
XFILL_10_DFFSR_18 gnd vdd FILL
XFILL_10_DFFSR_29 gnd vdd FILL
XFILL_58_DFFSR_116 gnd vdd FILL
XFILL_58_DFFSR_127 gnd vdd FILL
XFILL_58_DFFSR_138 gnd vdd FILL
XFILL_67_DFFSR_5 gnd vdd FILL
XFILL_58_DFFSR_149 gnd vdd FILL
XFILL_50_DFFSR_17 gnd vdd FILL
XFILL_1_DFFSR_109 gnd vdd FILL
XFILL_50_DFFSR_28 gnd vdd FILL
XFILL_50_DFFSR_39 gnd vdd FILL
XFILL_8_5_2 gnd vdd FILL
XFILL_7_0_1 gnd vdd FILL
XFILL_12_DFFSR_250 gnd vdd FILL
XFILL_12_DFFSR_261 gnd vdd FILL
XFILL_5_DFFSR_108 gnd vdd FILL
XFILL_12_DFFSR_272 gnd vdd FILL
XFILL_25_CLKBUF1_11 gnd vdd FILL
XFILL_5_DFFSR_119 gnd vdd FILL
XFILL_7_MUX2X1_9 gnd vdd FILL
XFILL_25_CLKBUF1_22 gnd vdd FILL
XFILL_25_CLKBUF1_33 gnd vdd FILL
XFILL_0_AOI21X1_4 gnd vdd FILL
XFILL_10_BUFX4_70 gnd vdd FILL
XFILL_16_DFFSR_260 gnd vdd FILL
XFILL_9_DFFSR_107 gnd vdd FILL
XFILL_16_DFFSR_271 gnd vdd FILL
XFILL_10_BUFX4_81 gnd vdd FILL
XFILL_8_CLKBUF1_15 gnd vdd FILL
XFILL_10_BUFX4_92 gnd vdd FILL
XFILL_13_MUX2X1_16 gnd vdd FILL
XFILL_9_DFFSR_118 gnd vdd FILL
XFILL_8_CLKBUF1_26 gnd vdd FILL
XFILL_44_7_0 gnd vdd FILL
XFILL_8_CLKBUF1_37 gnd vdd FILL
XFILL_9_DFFSR_129 gnd vdd FILL
XFILL_13_MUX2X1_27 gnd vdd FILL
XFILL_3_AOI21X1_12 gnd vdd FILL
XFILL_16_4_2 gnd vdd FILL
XFILL_13_MUX2X1_38 gnd vdd FILL
XFILL_4_AOI21X1_3 gnd vdd FILL
XFILL_13_MUX2X1_49 gnd vdd FILL
XFILL_3_AOI21X1_23 gnd vdd FILL
XFILL_3_AOI21X1_34 gnd vdd FILL
XFILL_43_DFFSR_160 gnd vdd FILL
XFILL_3_AOI21X1_45 gnd vdd FILL
XFILL_13_OAI22X1_14 gnd vdd FILL
XFILL_3_AOI21X1_56 gnd vdd FILL
XFILL_3_AOI21X1_67 gnd vdd FILL
XOAI21X1_15 INVX1_208/Y OAI21X1_5/B OAI21X1_15/C gnd NOR2X1_77/A vdd OAI21X1
XFILL_43_DFFSR_171 gnd vdd FILL
XFILL_3_AOI21X1_78 gnd vdd FILL
XOAI21X1_26 INVX1_190/Y OAI21X1_7/B NAND3X1_3/Y gnd NOR2X1_95/A vdd OAI21X1
XFILL_13_OAI22X1_25 gnd vdd FILL
XFILL_17_MUX2X1_15 gnd vdd FILL
XFILL_43_DFFSR_182 gnd vdd FILL
XFILL_43_DFFSR_193 gnd vdd FILL
XOAI21X1_37 INVX1_139/Y OAI21X1_37/B AND2X2_8/B gnd OAI21X1_38/C vdd OAI21X1
XFILL_13_OAI22X1_36 gnd vdd FILL
XFILL_13_OAI22X1_47 gnd vdd FILL
XOAI21X1_48 OAI21X1_48/A OAI21X1_48/B AOI22X1_1/C gnd NOR2X1_45/B vdd OAI21X1
XFILL_6_NOR2X1_100 gnd vdd FILL
XFILL_17_MUX2X1_26 gnd vdd FILL
XFILL_17_MUX2X1_37 gnd vdd FILL
XFILL_6_NOR2X1_111 gnd vdd FILL
XFILL_8_AOI21X1_2 gnd vdd FILL
XFILL_17_MUX2X1_48 gnd vdd FILL
XFILL_6_NOR2X1_122 gnd vdd FILL
XFILL_17_MUX2X1_59 gnd vdd FILL
XFILL_6_NOR2X1_133 gnd vdd FILL
XFILL_2_DFFSR_17 gnd vdd FILL
XFILL_13_NAND3X1_102 gnd vdd FILL
XFILL_6_NOR2X1_144 gnd vdd FILL
XFILL_2_DFFSR_28 gnd vdd FILL
XFILL_47_DFFSR_170 gnd vdd FILL
XFILL_13_NAND3X1_113 gnd vdd FILL
XFILL_6_NOR2X1_155 gnd vdd FILL
XFILL_5_NOR3X1_19 gnd vdd FILL
XFILL_6_INVX1_4 gnd vdd FILL
XFILL_6_NOR2X1_166 gnd vdd FILL
XFILL_2_DFFSR_39 gnd vdd FILL
XFILL_13_NAND3X1_124 gnd vdd FILL
XFILL_47_DFFSR_181 gnd vdd FILL
XFILL_21_DFFSR_106 gnd vdd FILL
XFILL_6_NOR2X1_177 gnd vdd FILL
XFILL_47_DFFSR_192 gnd vdd FILL
XFILL_6_NOR2X1_188 gnd vdd FILL
XFILL_6_NOR2X1_199 gnd vdd FILL
XFILL_21_DFFSR_117 gnd vdd FILL
XFILL_21_DFFSR_128 gnd vdd FILL
XFILL_12_NAND3X1_90 gnd vdd FILL
XFILL_4_INVX1_60 gnd vdd FILL
XFILL_21_DFFSR_139 gnd vdd FILL
XFILL_10_NOR2X1_205 gnd vdd FILL
XFILL_4_INVX1_71 gnd vdd FILL
XFILL_4_INVX1_82 gnd vdd FILL
XFILL_4_INVX1_93 gnd vdd FILL
XFILL_9_NOR3X1_18 gnd vdd FILL
XFILL_9_NOR3X1_29 gnd vdd FILL
XFILL_25_DFFSR_105 gnd vdd FILL
XFILL_25_DFFSR_116 gnd vdd FILL
XFILL_23_MUX2X1_102 gnd vdd FILL
XFILL_11_MUX2X1_3 gnd vdd FILL
XFILL_23_MUX2X1_113 gnd vdd FILL
XFILL_25_DFFSR_127 gnd vdd FILL
XFILL_25_DFFSR_138 gnd vdd FILL
XFILL_25_DFFSR_149 gnd vdd FILL
XFILL_23_MUX2X1_124 gnd vdd FILL
XFILL_4_NAND3X1_107 gnd vdd FILL
XFILL_23_MUX2X1_135 gnd vdd FILL
XFILL_23_MUX2X1_146 gnd vdd FILL
XFILL_4_NAND3X1_118 gnd vdd FILL
XFILL_23_MUX2X1_157 gnd vdd FILL
XFILL_4_NAND3X1_129 gnd vdd FILL
XFILL_23_MUX2X1_168 gnd vdd FILL
XFILL_29_DFFSR_104 gnd vdd FILL
XFILL_6_MUX2X1_106 gnd vdd FILL
XFILL_6_MUX2X1_117 gnd vdd FILL
XFILL_29_DFFSR_115 gnd vdd FILL
XFILL_23_MUX2X1_179 gnd vdd FILL
XFILL_6_MUX2X1_128 gnd vdd FILL
XFILL_29_DFFSR_126 gnd vdd FILL
XFILL_6_MUX2X1_139 gnd vdd FILL
XFILL_29_DFFSR_137 gnd vdd FILL
XFILL_2_BUFX4_80 gnd vdd FILL
XFILL_19_DFFSR_40 gnd vdd FILL
XFILL_19_DFFSR_51 gnd vdd FILL
XFILL_29_DFFSR_148 gnd vdd FILL
XFILL_2_BUFX4_91 gnd vdd FILL
XFILL_19_DFFSR_62 gnd vdd FILL
XFILL_3_OAI22X1_20 gnd vdd FILL
XFILL_29_DFFSR_159 gnd vdd FILL
XFILL_3_OAI22X1_31 gnd vdd FILL
XFILL_19_DFFSR_73 gnd vdd FILL
XFILL_66_3_2 gnd vdd FILL
XFILL_19_DFFSR_84 gnd vdd FILL
XFILL_3_OAI22X1_42 gnd vdd FILL
XFILL_21_NOR3X1_17 gnd vdd FILL
XFILL_7_OAI21X1_11 gnd vdd FILL
XFILL_19_DFFSR_95 gnd vdd FILL
XFILL_21_NOR3X1_28 gnd vdd FILL
XFILL_21_NOR3X1_39 gnd vdd FILL
XFILL_7_OAI21X1_22 gnd vdd FILL
XFILL_71_DFFSR_206 gnd vdd FILL
XFILL_7_OAI21X1_33 gnd vdd FILL
XFILL_71_DFFSR_217 gnd vdd FILL
XFILL_7_OAI21X1_44 gnd vdd FILL
XFILL_71_DFFSR_228 gnd vdd FILL
XFILL_59_DFFSR_50 gnd vdd FILL
XFILL_20_MUX2X1_1 gnd vdd FILL
XFILL_59_DFFSR_61 gnd vdd FILL
XFILL_35_7_0 gnd vdd FILL
XFILL_71_DFFSR_239 gnd vdd FILL
XFILL_59_DFFSR_72 gnd vdd FILL
XFILL_59_DFFSR_83 gnd vdd FILL
XFILL_25_NOR3X1_16 gnd vdd FILL
XFILL_25_NOR3X1_27 gnd vdd FILL
XFILL_59_DFFSR_94 gnd vdd FILL
XFILL_25_NOR3X1_38 gnd vdd FILL
XFILL_25_NOR3X1_49 gnd vdd FILL
XFILL_75_DFFSR_205 gnd vdd FILL
XFILL_0_NOR2X1_200 gnd vdd FILL
XFILL_75_DFFSR_216 gnd vdd FILL
XFILL_4_NOR2X1_4 gnd vdd FILL
XFILL_75_DFFSR_227 gnd vdd FILL
XFILL_10_DFFSR_160 gnd vdd FILL
XFILL_75_DFFSR_238 gnd vdd FILL
XFILL_75_DFFSR_249 gnd vdd FILL
XFILL_29_NOR3X1_15 gnd vdd FILL
XFILL_10_DFFSR_171 gnd vdd FILL
XFILL_29_NOR3X1_26 gnd vdd FILL
XFILL_10_DFFSR_182 gnd vdd FILL
XFILL_10_DFFSR_193 gnd vdd FILL
XFILL_28_DFFSR_60 gnd vdd FILL
XFILL_29_NOR3X1_37 gnd vdd FILL
XFILL_29_NOR3X1_48 gnd vdd FILL
XFILL_28_DFFSR_71 gnd vdd FILL
XFILL_28_DFFSR_82 gnd vdd FILL
XFILL_79_DFFSR_204 gnd vdd FILL
XFILL_79_DFFSR_215 gnd vdd FILL
XFILL_28_DFFSR_93 gnd vdd FILL
XFILL_79_DFFSR_226 gnd vdd FILL
XFILL_14_CLKBUF1_40 gnd vdd FILL
XFILL_79_DFFSR_237 gnd vdd FILL
XFILL_14_DFFSR_170 gnd vdd FILL
XFILL_3_MUX2X1_2 gnd vdd FILL
XFILL_79_DFFSR_248 gnd vdd FILL
XFILL_3_CLKBUF1_2 gnd vdd FILL
XFILL_79_DFFSR_259 gnd vdd FILL
XFILL_14_DFFSR_181 gnd vdd FILL
XFILL_14_DFFSR_192 gnd vdd FILL
XFILL_68_DFFSR_70 gnd vdd FILL
XFILL_11_DFFSR_4 gnd vdd FILL
XFILL_68_DFFSR_81 gnd vdd FILL
XFILL_68_DFFSR_92 gnd vdd FILL
XFILL_7_CLKBUF1_1 gnd vdd FILL
XFILL_18_DFFSR_180 gnd vdd FILL
XFILL_49_DFFSR_2 gnd vdd FILL
XFILL_18_DFFSR_191 gnd vdd FILL
XFILL_0_NOR3X1_8 gnd vdd FILL
XFILL_37_DFFSR_80 gnd vdd FILL
XFILL_37_DFFSR_91 gnd vdd FILL
XFILL_60_DFFSR_260 gnd vdd FILL
XFILL_60_DFFSR_271 gnd vdd FILL
XFILL_57_3_2 gnd vdd FILL
XFILL_77_DFFSR_90 gnd vdd FILL
XFILL_33_DFFSR_8 gnd vdd FILL
XFILL_64_DFFSR_270 gnd vdd FILL
XFILL_26_7_0 gnd vdd FILL
XFILL_1_7_0 gnd vdd FILL
XFILL_12_MUX2X1_120 gnd vdd FILL
XFILL_0_OAI21X1_7 gnd vdd FILL
XFILL_12_MUX2X1_131 gnd vdd FILL
XFILL_12_MUX2X1_142 gnd vdd FILL
XFILL_12_MUX2X1_153 gnd vdd FILL
XFILL_12_MUX2X1_164 gnd vdd FILL
XFILL_12_MUX2X1_175 gnd vdd FILL
XFILL_12_MUX2X1_186 gnd vdd FILL
XFILL_42_DFFSR_205 gnd vdd FILL
XFILL_1_NOR2X1_20 gnd vdd FILL
XFILL_40_2_2 gnd vdd FILL
XFILL_42_DFFSR_216 gnd vdd FILL
XFILL_4_OAI21X1_6 gnd vdd FILL
XFILL_1_NOR2X1_31 gnd vdd FILL
XFILL_42_DFFSR_227 gnd vdd FILL
XFILL_1_NOR2X1_42 gnd vdd FILL
XFILL_1_NOR2X1_53 gnd vdd FILL
XFILL_42_DFFSR_238 gnd vdd FILL
XFILL_42_DFFSR_249 gnd vdd FILL
XFILL_1_NOR2X1_64 gnd vdd FILL
XFILL_1_NOR2X1_75 gnd vdd FILL
XFILL_1_NOR2X1_86 gnd vdd FILL
XFILL_1_NOR2X1_97 gnd vdd FILL
XFILL_46_DFFSR_204 gnd vdd FILL
XFILL_46_DFFSR_215 gnd vdd FILL
XFILL_5_NOR2X1_30 gnd vdd FILL
XFILL_8_OAI21X1_5 gnd vdd FILL
XFILL_46_DFFSR_226 gnd vdd FILL
XFILL_5_NOR2X1_41 gnd vdd FILL
XFILL_46_DFFSR_237 gnd vdd FILL
XFILL_5_NOR2X1_52 gnd vdd FILL
XFILL_46_DFFSR_248 gnd vdd FILL
XFILL_5_NOR2X1_63 gnd vdd FILL
XFILL_5_NOR2X1_74 gnd vdd FILL
XFILL_46_DFFSR_259 gnd vdd FILL
XFILL_5_NOR2X1_85 gnd vdd FILL
XFILL_73_DFFSR_104 gnd vdd FILL
XFILL_5_NOR2X1_96 gnd vdd FILL
XFILL_73_DFFSR_115 gnd vdd FILL
XFILL_73_DFFSR_126 gnd vdd FILL
XFILL_9_NOR2X1_40 gnd vdd FILL
XFILL_73_DFFSR_137 gnd vdd FILL
XFILL_13_OAI22X1_2 gnd vdd FILL
XFILL_73_DFFSR_148 gnd vdd FILL
XFILL_9_NOR2X1_51 gnd vdd FILL
XFILL_9_NOR2X1_62 gnd vdd FILL
XFILL_73_DFFSR_159 gnd vdd FILL
XFILL_9_NOR2X1_73 gnd vdd FILL
XFILL_9_NOR2X1_84 gnd vdd FILL
XFILL_9_NOR2X1_95 gnd vdd FILL
XFILL_77_DFFSR_103 gnd vdd FILL
XFILL_6_8 gnd vdd FILL
XFILL_77_DFFSR_114 gnd vdd FILL
XFILL_77_DFFSR_125 gnd vdd FILL
XFILL_77_DFFSR_136 gnd vdd FILL
XFILL_15_NAND3X1_12 gnd vdd FILL
XFILL_17_OAI22X1_1 gnd vdd FILL
XFILL_77_DFFSR_147 gnd vdd FILL
XFILL_77_DFFSR_158 gnd vdd FILL
XFILL_2_MUX2X1_170 gnd vdd FILL
XFILL_15_NAND3X1_23 gnd vdd FILL
XFILL_48_3_2 gnd vdd FILL
XFILL_77_DFFSR_169 gnd vdd FILL
XFILL_15_NAND3X1_34 gnd vdd FILL
XFILL_2_MUX2X1_181 gnd vdd FILL
XFILL_2_MUX2X1_192 gnd vdd FILL
XFILL_15_NAND3X1_45 gnd vdd FILL
XFILL_15_NAND3X1_56 gnd vdd FILL
XFILL_35_CLKBUF1_12 gnd vdd FILL
XFILL_15_NAND3X1_67 gnd vdd FILL
XFILL_35_CLKBUF1_23 gnd vdd FILL
XFILL_15_NAND3X1_78 gnd vdd FILL
XFILL_15_NAND3X1_89 gnd vdd FILL
XFILL_35_CLKBUF1_34 gnd vdd FILL
XFILL_17_7_0 gnd vdd FILL
XFILL_31_DFFSR_270 gnd vdd FILL
XFILL_1_NAND2X1_8 gnd vdd FILL
XFILL_11_BUFX4_15 gnd vdd FILL
XFILL_11_BUFX4_26 gnd vdd FILL
XFILL_31_2_2 gnd vdd FILL
XFILL_11_BUFX4_37 gnd vdd FILL
XFILL_11_BUFX4_48 gnd vdd FILL
XFILL_5_NAND2X1_7 gnd vdd FILL
XFILL_11_BUFX4_59 gnd vdd FILL
XFILL_1_MUX2X1_60 gnd vdd FILL
XFILL_1_MUX2X1_71 gnd vdd FILL
XFILL_6_OAI22X1_19 gnd vdd FILL
XFILL_14_NAND3X1_103 gnd vdd FILL
XFILL_1_MUX2X1_82 gnd vdd FILL
XFILL_1_MUX2X1_93 gnd vdd FILL
XFILL_14_NAND3X1_114 gnd vdd FILL
XFILL_14_NAND3X1_125 gnd vdd FILL
XFILL_62_DFFSR_180 gnd vdd FILL
XDFFSR_18 DFFSR_18/Q DFFSR_88/CLK DFFSR_4/R vdd DFFSR_18/D gnd vdd DFFSR
XFILL_9_NAND2X1_6 gnd vdd FILL
XDFFSR_29 DFFSR_29/Q DFFSR_87/CLK DFFSR_87/R vdd DFFSR_29/D gnd vdd DFFSR
XFILL_62_DFFSR_191 gnd vdd FILL
XFILL_13_DFFSR_204 gnd vdd FILL
XFILL_13_DFFSR_215 gnd vdd FILL
XFILL_10_NAND3X1_4 gnd vdd FILL
XFILL_13_DFFSR_226 gnd vdd FILL
XFILL_5_MUX2X1_70 gnd vdd FILL
XFILL_5_MUX2X1_81 gnd vdd FILL
XFILL_13_DFFSR_237 gnd vdd FILL
XFILL_5_NAND3X1_40 gnd vdd FILL
XFILL_13_DFFSR_248 gnd vdd FILL
XFILL_5_NAND3X1_51 gnd vdd FILL
XFILL_5_NAND3X1_62 gnd vdd FILL
XFILL_5_MUX2X1_92 gnd vdd FILL
XFILL_50_DFFSR_2 gnd vdd FILL
XFILL_13_DFFSR_259 gnd vdd FILL
XFILL_9_NAND2X1_20 gnd vdd FILL
XFILL_5_NAND3X1_73 gnd vdd FILL
XFILL_9_NAND2X1_31 gnd vdd FILL
XFILL_40_DFFSR_104 gnd vdd FILL
XFILL_5_NAND3X1_84 gnd vdd FILL
XFILL_66_DFFSR_190 gnd vdd FILL
XFILL_9_NAND2X1_42 gnd vdd FILL
XFILL_14_NAND3X1_3 gnd vdd FILL
XFILL_5_NAND3X1_95 gnd vdd FILL
XFILL_17_DFFSR_203 gnd vdd FILL
XFILL_9_NAND2X1_53 gnd vdd FILL
XFILL_40_DFFSR_115 gnd vdd FILL
XFILL_17_DFFSR_214 gnd vdd FILL
XFILL_40_DFFSR_126 gnd vdd FILL
XFILL_17_DFFSR_225 gnd vdd FILL
XFILL_9_NAND2X1_64 gnd vdd FILL
XFILL_40_DFFSR_137 gnd vdd FILL
XFILL_17_DFFSR_236 gnd vdd FILL
XFILL_5_INVX1_16 gnd vdd FILL
XFILL_9_NAND2X1_75 gnd vdd FILL
XFILL_9_MUX2X1_80 gnd vdd FILL
XFILL_40_DFFSR_148 gnd vdd FILL
XFILL_9_NAND2X1_86 gnd vdd FILL
XFILL_5_INVX1_27 gnd vdd FILL
XFILL_22_13 gnd vdd FILL
XFILL_9_MUX2X1_91 gnd vdd FILL
XCLKBUF1_16 BUFX4_4/Y gnd DFFSR_1/CLK vdd CLKBUF1
XFILL_5_NAND3X1_108 gnd vdd FILL
XFILL_17_DFFSR_247 gnd vdd FILL
XFILL_40_DFFSR_159 gnd vdd FILL
XFILL_5_INVX1_38 gnd vdd FILL
XFILL_17_DFFSR_258 gnd vdd FILL
XFILL_5_NAND3X1_119 gnd vdd FILL
XCLKBUF1_27 BUFX4_73/Y gnd DFFSR_76/CLK vdd CLKBUF1
XFILL_17_DFFSR_269 gnd vdd FILL
XFILL_6_AND2X2_8 gnd vdd FILL
XFILL_5_INVX1_49 gnd vdd FILL
XCLKBUF1_38 BUFX4_10/Y gnd DFFSR_58/CLK vdd CLKBUF1
XFILL_44_DFFSR_103 gnd vdd FILL
XFILL_44_DFFSR_114 gnd vdd FILL
XFILL_17_CLKBUF1_17 gnd vdd FILL
XFILL_17_CLKBUF1_28 gnd vdd FILL
XFILL_39_3_2 gnd vdd FILL
XFILL_44_DFFSR_125 gnd vdd FILL
XFILL_44_DFFSR_136 gnd vdd FILL
XFILL_17_CLKBUF1_39 gnd vdd FILL
XFILL_12_AOI21X1_14 gnd vdd FILL
XFILL_44_DFFSR_147 gnd vdd FILL
XFILL_44_DFFSR_158 gnd vdd FILL
XBUFX4_70 INVX8_2/Y gnd MUX2X1_6/B vdd BUFX4
XFILL_12_AOI21X1_25 gnd vdd FILL
XFILL_44_DFFSR_169 gnd vdd FILL
XBUFX4_81 INVX8_4/Y gnd BUFX4_81/Y vdd BUFX4
XFILL_12_AOI21X1_36 gnd vdd FILL
XBUFX4_92 BUFX4_92/A gnd BUFX4_92/Y vdd BUFX4
XFILL_12_AOI21X1_47 gnd vdd FILL
XFILL_2_DFFSR_7 gnd vdd FILL
XFILL_48_DFFSR_102 gnd vdd FILL
XFILL_12_AOI21X1_58 gnd vdd FILL
XFILL_15_DFFSR_5 gnd vdd FILL
XFILL_12_AOI21X1_69 gnd vdd FILL
XFILL_48_DFFSR_113 gnd vdd FILL
XFILL_48_DFFSR_124 gnd vdd FILL
XFILL_3_BUFX4_14 gnd vdd FILL
XFILL_48_DFFSR_135 gnd vdd FILL
XFILL_72_DFFSR_6 gnd vdd FILL
XFILL_3_BUFX4_25 gnd vdd FILL
XFILL_48_DFFSR_146 gnd vdd FILL
XFILL_3_BUFX4_36 gnd vdd FILL
XFILL_48_DFFSR_157 gnd vdd FILL
XFILL_3_BUFX4_47 gnd vdd FILL
XFILL_10_AOI22X1_9 gnd vdd FILL
XFILL_48_DFFSR_168 gnd vdd FILL
XFILL_3_BUFX4_58 gnd vdd FILL
XFILL_48_DFFSR_179 gnd vdd FILL
XFILL_3_BUFX4_69 gnd vdd FILL
XFILL_21_MUX2X1_90 gnd vdd FILL
XFILL_50_5_0 gnd vdd FILL
XFILL_22_2_2 gnd vdd FILL
XFILL_14_AOI22X1_8 gnd vdd FILL
XFILL_24_CLKBUF1_30 gnd vdd FILL
XFILL_24_CLKBUF1_41 gnd vdd FILL
XFILL_0_NAND3X1_104 gnd vdd FILL
XFILL_0_NAND3X1_115 gnd vdd FILL
XFILL_18_AOI22X1_7 gnd vdd FILL
XFILL_37_DFFSR_9 gnd vdd FILL
XFILL_0_NAND3X1_126 gnd vdd FILL
XFILL_7_CLKBUF1_12 gnd vdd FILL
XFILL_7_CLKBUF1_23 gnd vdd FILL
XFILL_10_AND2X2_2 gnd vdd FILL
XFILL_7_CLKBUF1_34 gnd vdd FILL
XFILL_29_DFFSR_16 gnd vdd FILL
XFILL_29_DFFSR_27 gnd vdd FILL
XFILL_15_MUX2X1_108 gnd vdd FILL
XFILL_15_MUX2X1_119 gnd vdd FILL
XFILL_2_AOI21X1_20 gnd vdd FILL
XFILL_29_DFFSR_38 gnd vdd FILL
XFILL_2_AOI21X1_31 gnd vdd FILL
XFILL_29_DFFSR_49 gnd vdd FILL
XFILL_2_AOI21X1_42 gnd vdd FILL
XFILL_12_OAI22X1_11 gnd vdd FILL
XFILL_2_AOI21X1_53 gnd vdd FILL
XFILL_12_OAI22X1_22 gnd vdd FILL
XFILL_2_AOI21X1_64 gnd vdd FILL
XFILL_2_AOI21X1_75 gnd vdd FILL
XFILL_33_DFFSR_190 gnd vdd FILL
XFILL_12_OAI22X1_33 gnd vdd FILL
XFILL_69_DFFSR_15 gnd vdd FILL
XFILL_12_OAI22X1_44 gnd vdd FILL
XFILL_69_DFFSR_26 gnd vdd FILL
XFILL_69_DFFSR_37 gnd vdd FILL
XFILL_69_DFFSR_48 gnd vdd FILL
XFILL_5_NOR2X1_130 gnd vdd FILL
XFILL_69_DFFSR_59 gnd vdd FILL
XFILL_5_NOR2X1_141 gnd vdd FILL
XFILL_58_6_0 gnd vdd FILL
XFILL_5_NOR2X1_152 gnd vdd FILL
XFILL_5_NOR2X1_163 gnd vdd FILL
XFILL_5_NOR2X1_174 gnd vdd FILL
XFILL_5_3_2 gnd vdd FILL
XFILL_11_DFFSR_103 gnd vdd FILL
XFILL_11_DFFSR_114 gnd vdd FILL
XFILL_5_NOR2X1_185 gnd vdd FILL
XFILL_5_NOR2X1_196 gnd vdd FILL
XFILL_11_DFFSR_125 gnd vdd FILL
XFILL_11_DFFSR_136 gnd vdd FILL
XFILL_38_DFFSR_14 gnd vdd FILL
XFILL_11_DFFSR_147 gnd vdd FILL
XFILL_11_DFFSR_158 gnd vdd FILL
XFILL_38_DFFSR_25 gnd vdd FILL
XFILL_38_DFFSR_36 gnd vdd FILL
XFILL_11_DFFSR_169 gnd vdd FILL
XFILL_38_DFFSR_47 gnd vdd FILL
XFILL_15_DFFSR_102 gnd vdd FILL
XFILL_38_DFFSR_58 gnd vdd FILL
XFILL_38_DFFSR_69 gnd vdd FILL
XFILL_15_DFFSR_113 gnd vdd FILL
XFILL_15_DFFSR_124 gnd vdd FILL
XFILL_22_MUX2X1_110 gnd vdd FILL
XFILL_22_MUX2X1_121 gnd vdd FILL
XFILL_15_DFFSR_135 gnd vdd FILL
XFILL_15_DFFSR_146 gnd vdd FILL
XFILL_78_DFFSR_13 gnd vdd FILL
XFILL_15_DFFSR_157 gnd vdd FILL
XFILL_78_DFFSR_24 gnd vdd FILL
XFILL_22_MUX2X1_132 gnd vdd FILL
XFILL_78_DFFSR_35 gnd vdd FILL
XFILL_41_5_0 gnd vdd FILL
XFILL_15_DFFSR_168 gnd vdd FILL
XFILL_22_MUX2X1_143 gnd vdd FILL
XFILL_78_DFFSR_46 gnd vdd FILL
XFILL_22_MUX2X1_154 gnd vdd FILL
XFILL_13_2_2 gnd vdd FILL
XFILL_22_MUX2X1_165 gnd vdd FILL
XFILL_15_DFFSR_179 gnd vdd FILL
XFILL_78_DFFSR_57 gnd vdd FILL
XFILL_5_MUX2X1_103 gnd vdd FILL
XFILL_19_DFFSR_101 gnd vdd FILL
XFILL_22_MUX2X1_176 gnd vdd FILL
XFILL_5_MUX2X1_114 gnd vdd FILL
XFILL_78_DFFSR_68 gnd vdd FILL
XFILL_19_DFFSR_112 gnd vdd FILL
XFILL_5_MUX2X1_125 gnd vdd FILL
XFILL_22_MUX2X1_187 gnd vdd FILL
XFILL_78_DFFSR_79 gnd vdd FILL
XFILL_19_DFFSR_123 gnd vdd FILL
XINVX1_2 INVX1_2/A gnd INVX1_2/Y vdd INVX1
XFILL_5_MUX2X1_136 gnd vdd FILL
XFILL_1_INVX1_20 gnd vdd FILL
XFILL_19_DFFSR_134 gnd vdd FILL
XFILL_1_INVX1_31 gnd vdd FILL
XFILL_19_DFFSR_145 gnd vdd FILL
XFILL_1_INVX1_42 gnd vdd FILL
XFILL_5_MUX2X1_147 gnd vdd FILL
XFILL_19_DFFSR_156 gnd vdd FILL
XFILL_5_MUX2X1_158 gnd vdd FILL
XFILL_2_AND2X2_1 gnd vdd FILL
XFILL_19_DFFSR_167 gnd vdd FILL
XFILL_1_INVX1_53 gnd vdd FILL
XFILL_5_MUX2X1_169 gnd vdd FILL
XFILL_19_DFFSR_178 gnd vdd FILL
XFILL_1_INVX1_64 gnd vdd FILL
XFILL_11_NOR3X1_14 gnd vdd FILL
XFILL_47_DFFSR_12 gnd vdd FILL
XFILL_1_INVX1_75 gnd vdd FILL
XFILL_1_INVX1_86 gnd vdd FILL
XFILL_2_OAI22X1_50 gnd vdd FILL
XFILL_19_DFFSR_189 gnd vdd FILL
XFILL_11_NOR3X1_25 gnd vdd FILL
XFILL_1_INVX1_97 gnd vdd FILL
XFILL_11_NOR3X1_36 gnd vdd FILL
XFILL_47_DFFSR_23 gnd vdd FILL
XFILL_47_DFFSR_34 gnd vdd FILL
XFILL_6_OAI21X1_30 gnd vdd FILL
XFILL_11_NOR3X1_47 gnd vdd FILL
XFILL_18_NOR3X1_9 gnd vdd FILL
XFILL_61_DFFSR_203 gnd vdd FILL
XFILL_47_DFFSR_45 gnd vdd FILL
XFILL_47_DFFSR_56 gnd vdd FILL
XFILL_6_OAI21X1_41 gnd vdd FILL
XFILL_61_DFFSR_214 gnd vdd FILL
XFILL_47_DFFSR_67 gnd vdd FILL
XFILL_61_DFFSR_225 gnd vdd FILL
XFILL_61_DFFSR_236 gnd vdd FILL
XFILL_4_BUFX4_105 gnd vdd FILL
XFILL_47_DFFSR_78 gnd vdd FILL
XFILL_47_DFFSR_89 gnd vdd FILL
XFILL_61_DFFSR_247 gnd vdd FILL
XFILL_15_NOR3X1_13 gnd vdd FILL
XFILL_87_DFFSR_11 gnd vdd FILL
XFILL_61_DFFSR_258 gnd vdd FILL
XFILL_61_DFFSR_269 gnd vdd FILL
XFILL_15_NOR3X1_24 gnd vdd FILL
XFILL_87_DFFSR_22 gnd vdd FILL
XFILL_15_NOR3X1_35 gnd vdd FILL
XFILL_15_NOR3X1_46 gnd vdd FILL
XFILL_87_DFFSR_33 gnd vdd FILL
XFILL_65_DFFSR_202 gnd vdd FILL
XFILL_87_DFFSR_44 gnd vdd FILL
XFILL_87_DFFSR_55 gnd vdd FILL
XFILL_65_DFFSR_213 gnd vdd FILL
XFILL_16_DFFSR_11 gnd vdd FILL
XFILL_16_DFFSR_22 gnd vdd FILL
XFILL_87_DFFSR_66 gnd vdd FILL
XFILL_65_DFFSR_224 gnd vdd FILL
XFILL_87_DFFSR_77 gnd vdd FILL
XFILL_65_DFFSR_235 gnd vdd FILL
XFILL_8_BUFX4_104 gnd vdd FILL
XFILL_16_DFFSR_33 gnd vdd FILL
XFILL_87_DFFSR_88 gnd vdd FILL
XFILL_65_DFFSR_246 gnd vdd FILL
XFILL_16_DFFSR_44 gnd vdd FILL
XFILL_16_DFFSR_55 gnd vdd FILL
XFILL_87_DFFSR_99 gnd vdd FILL
XFILL_4_5 gnd vdd FILL
XFILL_19_NOR3X1_12 gnd vdd FILL
XFILL_65_DFFSR_257 gnd vdd FILL
XFILL_65_DFFSR_268 gnd vdd FILL
XFILL_16_DFFSR_66 gnd vdd FILL
XFILL_19_NOR3X1_23 gnd vdd FILL
XFILL_12_INVX8_3 gnd vdd FILL
XFILL_19_NOR3X1_34 gnd vdd FILL
XFILL_16_DFFSR_77 gnd vdd FILL
XFILL_20_CLKBUF1_9 gnd vdd FILL
XFILL_69_DFFSR_201 gnd vdd FILL
XFILL_19_NOR3X1_45 gnd vdd FILL
XFILL_49_6_0 gnd vdd FILL
XFILL_16_DFFSR_88 gnd vdd FILL
XFILL_60_7 gnd vdd FILL
XFILL_16_DFFSR_99 gnd vdd FILL
XFILL_69_DFFSR_212 gnd vdd FILL
XFILL_56_DFFSR_10 gnd vdd FILL
XFILL_56_DFFSR_21 gnd vdd FILL
XFILL_69_DFFSR_223 gnd vdd FILL
XFILL_69_DFFSR_234 gnd vdd FILL
XFILL_56_DFFSR_32 gnd vdd FILL
XFILL_69_DFFSR_245 gnd vdd FILL
XFILL_27_NOR3X1_7 gnd vdd FILL
XFILL_56_DFFSR_43 gnd vdd FILL
XFILL_69_DFFSR_256 gnd vdd FILL
XFILL_56_DFFSR_54 gnd vdd FILL
XFILL_69_DFFSR_267 gnd vdd FILL
XFILL_56_DFFSR_65 gnd vdd FILL
XFILL_56_DFFSR_76 gnd vdd FILL
XFILL_24_CLKBUF1_8 gnd vdd FILL
XFILL_56_DFFSR_87 gnd vdd FILL
XFILL_2_NOR2X1_18 gnd vdd FILL
XFILL_56_DFFSR_98 gnd vdd FILL
XFILL_46_5 gnd vdd FILL
XFILL_63_1_2 gnd vdd FILL
XFILL_8_NAND3X1_17 gnd vdd FILL
XFILL_2_NOR2X1_29 gnd vdd FILL
XFILL_8_NAND3X1_28 gnd vdd FILL
XFILL_8_NAND3X1_39 gnd vdd FILL
XFILL_54_DFFSR_3 gnd vdd FILL
XFILL_1_NOR2X1_8 gnd vdd FILL
XFILL_25_DFFSR_20 gnd vdd FILL
XFILL_28_CLKBUF1_7 gnd vdd FILL
XFILL_25_DFFSR_31 gnd vdd FILL
XFILL_25_DFFSR_42 gnd vdd FILL
XFILL_6_NOR2X1_17 gnd vdd FILL
XFILL_6_NOR2X1_28 gnd vdd FILL
XFILL_25_DFFSR_53 gnd vdd FILL
XFILL_32_5_0 gnd vdd FILL
XFILL_25_DFFSR_64 gnd vdd FILL
XFILL_25_DFFSR_75 gnd vdd FILL
XFILL_6_NOR2X1_39 gnd vdd FILL
XFILL_25_DFFSR_86 gnd vdd FILL
XFILL_25_DFFSR_97 gnd vdd FILL
XFILL_65_DFFSR_30 gnd vdd FILL
XFILL_65_DFFSR_41 gnd vdd FILL
XFILL_0_MUX2X1_6 gnd vdd FILL
XFILL_65_DFFSR_52 gnd vdd FILL
XFILL_65_DFFSR_63 gnd vdd FILL
XFILL_65_DFFSR_74 gnd vdd FILL
XFILL_65_DFFSR_85 gnd vdd FILL
XFILL_65_DFFSR_96 gnd vdd FILL
XFILL_1_NAND2X1_19 gnd vdd FILL
XFILL_15_NAND3X1_104 gnd vdd FILL
XFILL_6_DFFSR_8 gnd vdd FILL
XFILL_15_NAND3X1_115 gnd vdd FILL
XFILL_15_NAND3X1_126 gnd vdd FILL
XFILL_8_DFFSR_10 gnd vdd FILL
XFILL_8_DFFSR_21 gnd vdd FILL
XFILL_19_DFFSR_6 gnd vdd FILL
XFILL_8_DFFSR_32 gnd vdd FILL
XFILL_8_DFFSR_43 gnd vdd FILL
XFILL_76_DFFSR_7 gnd vdd FILL
XFILL_8_DFFSR_54 gnd vdd FILL
XFILL_34_DFFSR_40 gnd vdd FILL
XFILL_8_DFFSR_65 gnd vdd FILL
XFILL_8_DFFSR_76 gnd vdd FILL
XFILL_34_DFFSR_51 gnd vdd FILL
XFILL_11_MUX2X1_150 gnd vdd FILL
XFILL_8_DFFSR_87 gnd vdd FILL
XFILL_34_DFFSR_62 gnd vdd FILL
XFILL_11_MUX2X1_161 gnd vdd FILL
XFILL_8_DFFSR_98 gnd vdd FILL
XFILL_34_DFFSR_73 gnd vdd FILL
XFILL_11_MUX2X1_172 gnd vdd FILL
XFILL_34_DFFSR_84 gnd vdd FILL
XFILL_34_DFFSR_95 gnd vdd FILL
XFILL_11_MUX2X1_183 gnd vdd FILL
XFILL_32_DFFSR_202 gnd vdd FILL
XFILL_11_MUX2X1_194 gnd vdd FILL
XFILL_32_DFFSR_213 gnd vdd FILL
XFILL_32_DFFSR_224 gnd vdd FILL
XFILL_32_DFFSR_235 gnd vdd FILL
XFILL_74_DFFSR_50 gnd vdd FILL
XFILL_32_DFFSR_246 gnd vdd FILL
XFILL_74_DFFSR_61 gnd vdd FILL
XFILL_6_NAND3X1_109 gnd vdd FILL
XFILL_1_DFFSR_270 gnd vdd FILL
XFILL_32_DFFSR_257 gnd vdd FILL
XFILL_74_DFFSR_72 gnd vdd FILL
XFILL_32_DFFSR_268 gnd vdd FILL
XFILL_74_DFFSR_83 gnd vdd FILL
XFILL_74_DFFSR_94 gnd vdd FILL
XFILL_36_DFFSR_201 gnd vdd FILL
XFILL_27_CLKBUF1_18 gnd vdd FILL
XFILL_27_CLKBUF1_29 gnd vdd FILL
XFILL_36_DFFSR_212 gnd vdd FILL
XFILL_36_DFFSR_223 gnd vdd FILL
XFILL_36_DFFSR_234 gnd vdd FILL
XFILL_36_DFFSR_245 gnd vdd FILL
XFILL_36_DFFSR_256 gnd vdd FILL
XFILL_54_1_2 gnd vdd FILL
XFILL_36_DFFSR_267 gnd vdd FILL
XFILL_14_NOR3X1_2 gnd vdd FILL
XFILL_2_MUX2X1_14 gnd vdd FILL
XFILL_2_MUX2X1_25 gnd vdd FILL
XFILL_63_DFFSR_101 gnd vdd FILL
XFILL_43_DFFSR_60 gnd vdd FILL
XFILL_2_MUX2X1_36 gnd vdd FILL
XFILL_63_DFFSR_112 gnd vdd FILL
XFILL_2_MUX2X1_47 gnd vdd FILL
XFILL_43_DFFSR_71 gnd vdd FILL
XFILL_63_DFFSR_123 gnd vdd FILL
XFILL_43_DFFSR_82 gnd vdd FILL
XFILL_5_AOI21X1_19 gnd vdd FILL
XFILL_2_MUX2X1_58 gnd vdd FILL
XFILL_63_DFFSR_134 gnd vdd FILL
XFILL_2_MUX2X1_69 gnd vdd FILL
XFILL_43_DFFSR_93 gnd vdd FILL
XFILL_63_DFFSR_145 gnd vdd FILL
XFILL_10_NAND3X1_100 gnd vdd FILL
XFILL_63_DFFSR_156 gnd vdd FILL
XFILL_10_NAND3X1_111 gnd vdd FILL
XFILL_63_DFFSR_167 gnd vdd FILL
XFILL_23_5_0 gnd vdd FILL
XFILL_10_NAND3X1_122 gnd vdd FILL
XFILL_6_MUX2X1_13 gnd vdd FILL
XFILL_63_DFFSR_178 gnd vdd FILL
XFILL_6_MUX2X1_24 gnd vdd FILL
XFILL_67_DFFSR_100 gnd vdd FILL
XFILL_63_DFFSR_189 gnd vdd FILL
XFILL_6_MUX2X1_35 gnd vdd FILL
XFILL_67_DFFSR_111 gnd vdd FILL
XFILL_8_NOR2X1_107 gnd vdd FILL
XFILL_83_DFFSR_70 gnd vdd FILL
XFILL_67_DFFSR_122 gnd vdd FILL
XFILL_6_MUX2X1_46 gnd vdd FILL
XFILL_8_NOR2X1_118 gnd vdd FILL
XFILL_67_DFFSR_133 gnd vdd FILL
XFILL_83_DFFSR_81 gnd vdd FILL
XFILL_6_MUX2X1_57 gnd vdd FILL
XFILL_83_DFFSR_92 gnd vdd FILL
XFILL_8_NOR2X1_129 gnd vdd FILL
XFILL_6_MUX2X1_68 gnd vdd FILL
XFILL_6_MUX2X1_79 gnd vdd FILL
XFILL_67_DFFSR_144 gnd vdd FILL
XFILL_10_OAI21X1_1 gnd vdd FILL
XFILL_14_NAND3X1_20 gnd vdd FILL
XFILL_67_DFFSR_155 gnd vdd FILL
XFILL_0_BUFX4_8 gnd vdd FILL
XFILL_12_DFFSR_70 gnd vdd FILL
XFILL_14_NAND3X1_31 gnd vdd FILL
XFILL_67_DFFSR_166 gnd vdd FILL
XFILL_67_DFFSR_177 gnd vdd FILL
XFILL_12_DFFSR_81 gnd vdd FILL
XFILL_14_NAND3X1_42 gnd vdd FILL
XFILL_13_BUFX4_6 gnd vdd FILL
XFILL_12_DFFSR_92 gnd vdd FILL
XFILL_14_NAND3X1_53 gnd vdd FILL
XFILL_67_DFFSR_188 gnd vdd FILL
XFILL_14_NAND3X1_64 gnd vdd FILL
XFILL_67_DFFSR_199 gnd vdd FILL
XFILL_34_CLKBUF1_20 gnd vdd FILL
XFILL_14_NAND3X1_75 gnd vdd FILL
XFILL_14_NAND3X1_86 gnd vdd FILL
XFILL_34_CLKBUF1_31 gnd vdd FILL
XFILL_14_NAND3X1_97 gnd vdd FILL
XFILL_34_CLKBUF1_42 gnd vdd FILL
XFILL_1_NAND3X1_105 gnd vdd FILL
XFILL_1_NAND3X1_116 gnd vdd FILL
XFILL_1_NAND3X1_127 gnd vdd FILL
XFILL_52_DFFSR_80 gnd vdd FILL
XFILL_52_DFFSR_91 gnd vdd FILL
XFILL_11_NOR2X1_80 gnd vdd FILL
XFILL_11_NOR2X1_91 gnd vdd FILL
XFILL_22_MUX2X1_11 gnd vdd FILL
XFILL_22_MUX2X1_22 gnd vdd FILL
XFILL_22_MUX2X1_33 gnd vdd FILL
XFILL_21_DFFSR_90 gnd vdd FILL
XFILL_6_6_0 gnd vdd FILL
XFILL_22_MUX2X1_44 gnd vdd FILL
XFILL_22_MUX2X1_55 gnd vdd FILL
XFILL_6_NOR3X1_1 gnd vdd FILL
XFILL_22_MUX2X1_66 gnd vdd FILL
XFILL_5_OAI22X1_16 gnd vdd FILL
XFILL_22_MUX2X1_77 gnd vdd FILL
XFILL_5_OAI22X1_27 gnd vdd FILL
XFILL_5_OAI22X1_38 gnd vdd FILL
XFILL_22_MUX2X1_88 gnd vdd FILL
XFILL_22_MUX2X1_99 gnd vdd FILL
XFILL_5_OAI22X1_49 gnd vdd FILL
XFILL_9_OAI21X1_18 gnd vdd FILL
XFILL_9_OAI21X1_29 gnd vdd FILL
XFILL_45_1_2 gnd vdd FILL
XFILL_4_NAND3X1_70 gnd vdd FILL
XFILL_30_DFFSR_101 gnd vdd FILL
XFILL_4_NAND3X1_81 gnd vdd FILL
XFILL_4_NAND3X1_92 gnd vdd FILL
XFILL_8_NAND2X1_50 gnd vdd FILL
XFILL_30_DFFSR_112 gnd vdd FILL
XFILL_14_5_0 gnd vdd FILL
XFILL_8_NAND2X1_61 gnd vdd FILL
XFILL_30_DFFSR_123 gnd vdd FILL
XFILL_4_DFFSR_80 gnd vdd FILL
XFILL_30_DFFSR_134 gnd vdd FILL
XFILL_8_NAND2X1_72 gnd vdd FILL
XFILL_30_DFFSR_145 gnd vdd FILL
XFILL_4_DFFSR_91 gnd vdd FILL
XFILL_8_NAND2X1_83 gnd vdd FILL
XFILL_30_DFFSR_156 gnd vdd FILL
XFILL_8_NAND2X1_94 gnd vdd FILL
XFILL_30_DFFSR_167 gnd vdd FILL
XFILL_16_INVX8_4 gnd vdd FILL
XFILL_30_DFFSR_178 gnd vdd FILL
XFILL_34_DFFSR_100 gnd vdd FILL
XFILL_30_DFFSR_189 gnd vdd FILL
XFILL_34_DFFSR_111 gnd vdd FILL
XFILL_16_CLKBUF1_14 gnd vdd FILL
XFILL_11_NAND2X1_2 gnd vdd FILL
XFILL_16_CLKBUF1_25 gnd vdd FILL
XFILL_34_DFFSR_122 gnd vdd FILL
XFILL_16_CLKBUF1_36 gnd vdd FILL
XFILL_34_DFFSR_133 gnd vdd FILL
XFILL_11_AOI21X1_11 gnd vdd FILL
XFILL_34_DFFSR_144 gnd vdd FILL
XFILL_34_DFFSR_155 gnd vdd FILL
XFILL_11_AOI21X1_22 gnd vdd FILL
XFILL_34_DFFSR_166 gnd vdd FILL
XFILL_34_DFFSR_177 gnd vdd FILL
XFILL_11_AOI21X1_33 gnd vdd FILL
XFILL_11_AOI21X1_44 gnd vdd FILL
XFILL_3_DFFSR_190 gnd vdd FILL
XAND2X2_2 AND2X2_2/A AND2X2_2/B gnd BUFX4_2/A vdd AND2X2
XFILL_34_DFFSR_188 gnd vdd FILL
XFILL_11_AOI21X1_55 gnd vdd FILL
XFILL_11_AOI21X1_66 gnd vdd FILL
XFILL_20_DFFSR_6 gnd vdd FILL
XFILL_38_DFFSR_110 gnd vdd FILL
XFILL_34_DFFSR_199 gnd vdd FILL
XFILL_11_AOI21X1_77 gnd vdd FILL
XFILL_38_DFFSR_121 gnd vdd FILL
XFILL_38_DFFSR_132 gnd vdd FILL
XFILL_38_DFFSR_143 gnd vdd FILL
XFILL_38_DFFSR_154 gnd vdd FILL
XFILL_58_DFFSR_4 gnd vdd FILL
XFILL_38_DFFSR_165 gnd vdd FILL
XFILL_38_DFFSR_176 gnd vdd FILL
XFILL_38_DFFSR_187 gnd vdd FILL
XFILL_30_NOR3X1_12 gnd vdd FILL
XFILL_30_NOR3X1_23 gnd vdd FILL
XFILL_30_NOR3X1_34 gnd vdd FILL
XFILL_38_DFFSR_198 gnd vdd FILL
XFILL_30_NOR3X1_45 gnd vdd FILL
XFILL_80_DFFSR_201 gnd vdd FILL
XFILL_80_DFFSR_212 gnd vdd FILL
XFILL_80_DFFSR_223 gnd vdd FILL
XFILL_2_2 gnd vdd FILL
XFILL_80_DFFSR_234 gnd vdd FILL
XFILL_80_DFFSR_245 gnd vdd FILL
XFILL_80_DFFSR_256 gnd vdd FILL
XFILL_80_DFFSR_267 gnd vdd FILL
XFILL_84_DFFSR_200 gnd vdd FILL
XFILL_84_DFFSR_211 gnd vdd FILL
XFILL_84_DFFSR_222 gnd vdd FILL
XFILL_11_AOI21X1_7 gnd vdd FILL
XFILL_0_BUFX4_18 gnd vdd FILL
XFILL_84_DFFSR_233 gnd vdd FILL
XFILL_84_DFFSR_244 gnd vdd FILL
XFILL_64_4_0 gnd vdd FILL
XFILL_0_BUFX4_29 gnd vdd FILL
XFILL_84_DFFSR_255 gnd vdd FILL
XFILL_6_CLKBUF1_20 gnd vdd FILL
XFILL_44_2 gnd vdd FILL
XFILL_36_1_2 gnd vdd FILL
XFILL_84_DFFSR_266 gnd vdd FILL
XFILL_6_CLKBUF1_31 gnd vdd FILL
XFILL_6_CLKBUF1_42 gnd vdd FILL
XFILL_14_MUX2X1_105 gnd vdd FILL
XFILL_14_MUX2X1_116 gnd vdd FILL
XFILL_0_INVX1_150 gnd vdd FILL
XFILL_14_MUX2X1_127 gnd vdd FILL
XFILL_0_INVX1_161 gnd vdd FILL
XFILL_15_AOI21X1_6 gnd vdd FILL
XFILL_1_AOI21X1_50 gnd vdd FILL
XFILL_14_MUX2X1_138 gnd vdd FILL
XFILL_0_INVX1_172 gnd vdd FILL
XFILL_14_MUX2X1_149 gnd vdd FILL
XFILL_0_INVX1_183 gnd vdd FILL
XFILL_1_AOI21X1_61 gnd vdd FILL
XFILL_1_AOI21X1_72 gnd vdd FILL
XFILL_11_OAI22X1_30 gnd vdd FILL
XFILL_0_INVX1_194 gnd vdd FILL
XFILL_11_OAI22X1_41 gnd vdd FILL
XFILL_15_OAI21X1_10 gnd vdd FILL
XFILL_15_OAI21X1_21 gnd vdd FILL
XFILL_4_INVX1_160 gnd vdd FILL
XFILL_15_OAI21X1_32 gnd vdd FILL
XFILL_4_INVX1_171 gnd vdd FILL
XFILL_15_OAI21X1_43 gnd vdd FILL
XFILL_4_INVX1_182 gnd vdd FILL
XFILL_4_NOR2X1_160 gnd vdd FILL
XFILL_4_INVX1_193 gnd vdd FILL
XFILL_4_NOR2X1_171 gnd vdd FILL
XFILL_4_NOR2X1_182 gnd vdd FILL
XFILL_4_NOR2X1_193 gnd vdd FILL
XFILL_66_DFFSR_19 gnd vdd FILL
XFILL_21_MUX2X1_140 gnd vdd FILL
XFILL_21_MUX2X1_151 gnd vdd FILL
XFILL_4_MUX2X1_100 gnd vdd FILL
XFILL_60_10 gnd vdd FILL
XFILL_21_MUX2X1_162 gnd vdd FILL
XFILL_21_MUX2X1_173 gnd vdd FILL
XFILL_4_MUX2X1_111 gnd vdd FILL
XFILL_21_MUX2X1_184 gnd vdd FILL
XFILL_4_MUX2X1_122 gnd vdd FILL
XNAND3X1_18 NAND3X1_18/A NAND3X1_18/B NOR2X1_103/Y gnd NOR3X1_44/B vdd NAND3X1
XNAND3X1_29 INVX1_136/Y OAI21X1_36/Y NAND3X1_29/C gnd AOI22X1_1/B vdd NAND3X1
XFILL_4_MUX2X1_133 gnd vdd FILL
XFILL_4_MUX2X1_144 gnd vdd FILL
XFILL_4_BUFX4_9 gnd vdd FILL
XFILL_4_MUX2X1_155 gnd vdd FILL
XFILL_4_MUX2X1_166 gnd vdd FILL
XFILL_4_MUX2X1_177 gnd vdd FILL
XFILL_4_MUX2X1_188 gnd vdd FILL
XFILL_35_DFFSR_18 gnd vdd FILL
XFILL_35_DFFSR_29 gnd vdd FILL
XNOR2X1_18 NOR2X1_18/A NOR2X1_19/B gnd NOR2X1_18/Y vdd NOR2X1
XNOR2X1_29 NOR3X1_52/C NOR2X1_37/B gnd NOR2X1_29/Y vdd NOR2X1
XFILL_51_DFFSR_200 gnd vdd FILL
XFILL_51_DFFSR_211 gnd vdd FILL
XFILL_55_4_0 gnd vdd FILL
XFILL_51_DFFSR_222 gnd vdd FILL
XFILL_27_1_2 gnd vdd FILL
XFILL_51_DFFSR_233 gnd vdd FILL
XFILL_2_1_2 gnd vdd FILL
XFILL_51_DFFSR_244 gnd vdd FILL
XFILL_51_DFFSR_255 gnd vdd FILL
XFILL_75_DFFSR_17 gnd vdd FILL
XFILL_75_DFFSR_28 gnd vdd FILL
XFILL_51_DFFSR_266 gnd vdd FILL
XFILL_75_DFFSR_39 gnd vdd FILL
XFILL_18_MUX2X1_7 gnd vdd FILL
XFILL_55_DFFSR_210 gnd vdd FILL
XFILL_55_DFFSR_221 gnd vdd FILL
XFILL_55_DFFSR_232 gnd vdd FILL
XFILL_55_DFFSR_243 gnd vdd FILL
XFILL_11_NAND3X1_101 gnd vdd FILL
XFILL_11_NAND3X1_112 gnd vdd FILL
XFILL_55_DFFSR_254 gnd vdd FILL
XFILL_11_NAND3X1_123 gnd vdd FILL
XFILL_55_DFFSR_265 gnd vdd FILL
XFILL_9_BUFX4_40 gnd vdd FILL
XFILL_10_CLKBUF1_6 gnd vdd FILL
XFILL_9_BUFX4_51 gnd vdd FILL
XFILL_44_DFFSR_16 gnd vdd FILL
XFILL_82_DFFSR_110 gnd vdd FILL
XFILL_9_BUFX4_62 gnd vdd FILL
XFILL_9_BUFX4_73 gnd vdd FILL
XFILL_82_DFFSR_121 gnd vdd FILL
XFILL_9_BUFX4_84 gnd vdd FILL
XFILL_0_BUFX2_5 gnd vdd FILL
XFILL_59_DFFSR_220 gnd vdd FILL
XFILL_10_0_2 gnd vdd FILL
XFILL_44_DFFSR_27 gnd vdd FILL
XFILL_82_DFFSR_132 gnd vdd FILL
XFILL_44_DFFSR_38 gnd vdd FILL
XFILL_59_DFFSR_231 gnd vdd FILL
XFILL_9_BUFX4_95 gnd vdd FILL
XFILL_82_DFFSR_143 gnd vdd FILL
XFILL_59_DFFSR_242 gnd vdd FILL
XFILL_44_DFFSR_49 gnd vdd FILL
XFILL_82_DFFSR_154 gnd vdd FILL
XFILL_59_DFFSR_253 gnd vdd FILL
XFILL_82_DFFSR_165 gnd vdd FILL
XFILL_59_DFFSR_264 gnd vdd FILL
XFILL_82_DFFSR_176 gnd vdd FILL
XFILL_59_DFFSR_275 gnd vdd FILL
XFILL_14_CLKBUF1_5 gnd vdd FILL
XFILL_2_DFFSR_202 gnd vdd FILL
XFILL_82_DFFSR_187 gnd vdd FILL
XFILL_2_DFFSR_213 gnd vdd FILL
XFILL_82_DFFSR_198 gnd vdd FILL
XFILL_84_DFFSR_15 gnd vdd FILL
XFILL_86_DFFSR_120 gnd vdd FILL
XFILL_7_NAND3X1_14 gnd vdd FILL
XFILL_84_DFFSR_26 gnd vdd FILL
XFILL_2_DFFSR_224 gnd vdd FILL
XFILL_86_DFFSR_131 gnd vdd FILL
XFILL_2_DFFSR_235 gnd vdd FILL
XFILL_7_NAND3X1_25 gnd vdd FILL
XFILL_84_DFFSR_37 gnd vdd FILL
XFILL_86_DFFSR_142 gnd vdd FILL
XFILL_84_DFFSR_48 gnd vdd FILL
XFILL_7_NAND3X1_36 gnd vdd FILL
XFILL_2_DFFSR_246 gnd vdd FILL
XFILL_2_NAND3X1_106 gnd vdd FILL
XFILL_86_DFFSR_153 gnd vdd FILL
XFILL_2_NAND3X1_117 gnd vdd FILL
XFILL_7_NAND3X1_47 gnd vdd FILL
XFILL_13_DFFSR_15 gnd vdd FILL
XFILL_2_DFFSR_257 gnd vdd FILL
XFILL_84_DFFSR_59 gnd vdd FILL
XFILL_10_BUFX4_100 gnd vdd FILL
XFILL_2_DFFSR_268 gnd vdd FILL
XFILL_2_NAND3X1_128 gnd vdd FILL
XFILL_7_NAND3X1_58 gnd vdd FILL
XFILL_13_DFFSR_26 gnd vdd FILL
XFILL_86_DFFSR_164 gnd vdd FILL
XFILL_7_NAND3X1_69 gnd vdd FILL
XFILL_86_DFFSR_175 gnd vdd FILL
XFILL_18_CLKBUF1_4 gnd vdd FILL
XFILL_6_DFFSR_201 gnd vdd FILL
XFILL_13_DFFSR_37 gnd vdd FILL
XFILL_86_DFFSR_186 gnd vdd FILL
XFILL_13_DFFSR_48 gnd vdd FILL
XFILL_3_NAND3X1_1 gnd vdd FILL
XFILL_86_DFFSR_197 gnd vdd FILL
XFILL_6_DFFSR_212 gnd vdd FILL
XFILL_13_DFFSR_59 gnd vdd FILL
XFILL_6_DFFSR_223 gnd vdd FILL
XFILL_6_DFFSR_234 gnd vdd FILL
XFILL_6_DFFSR_245 gnd vdd FILL
XFILL_53_DFFSR_14 gnd vdd FILL
XFILL_6_DFFSR_256 gnd vdd FILL
XFILL_6_DFFSR_267 gnd vdd FILL
XFILL_53_DFFSR_25 gnd vdd FILL
XFILL_53_DFFSR_36 gnd vdd FILL
XFILL_53_DFFSR_47 gnd vdd FILL
XFILL_53_DFFSR_58 gnd vdd FILL
XFILL_53_DFFSR_69 gnd vdd FILL
XMUX2X1_14 BUFX4_75/Y INVX1_27/Y MUX2X1_14/S gnd DFFSR_34/D vdd MUX2X1
XFILL_0_NAND2X1_16 gnd vdd FILL
XMUX2X1_25 BUFX4_71/Y INVX1_38/Y NOR2X1_9/B gnd MUX2X1_25/Y vdd MUX2X1
XFILL_0_NAND2X1_27 gnd vdd FILL
XFILL_46_4_0 gnd vdd FILL
XFILL_18_1_2 gnd vdd FILL
XMUX2X1_36 MUX2X1_7/B INVX1_49/Y NOR2X1_20/Y gnd MUX2X1_36/Y vdd MUX2X1
XFILL_0_NAND2X1_38 gnd vdd FILL
XMUX2X1_47 INVX1_60/Y MUX2X1_9/A NAND2X1_7/Y gnd MUX2X1_47/Y vdd MUX2X1
XNOR2X1_108 INVX2_3/A BUFX2_7/A gnd AND2X2_7/A vdd NOR2X1
XFILL_24_DFFSR_7 gnd vdd FILL
XFILL_22_DFFSR_13 gnd vdd FILL
XFILL_68_DFFSR_109 gnd vdd FILL
XFILL_0_NAND2X1_49 gnd vdd FILL
XNOR2X1_119 OAI21X1_39/B AOI22X1_3/A gnd OAI21X1_45/A vdd NOR2X1
XFILL_22_DFFSR_24 gnd vdd FILL
XFILL_81_DFFSR_8 gnd vdd FILL
XMUX2X1_58 INVX1_71/Y MUX2X1_66/A NAND2X1_9/Y gnd MUX2X1_58/Y vdd MUX2X1
XMUX2X1_69 INVX1_82/Y BUFX4_64/Y MUX2X1_71/S gnd MUX2X1_69/Y vdd MUX2X1
XFILL_22_DFFSR_35 gnd vdd FILL
XFILL_22_DFFSR_46 gnd vdd FILL
XFILL_22_DFFSR_57 gnd vdd FILL
XFILL_0_INVX2_5 gnd vdd FILL
XFILL_22_DFFSR_68 gnd vdd FILL
XFILL_22_DFFSR_79 gnd vdd FILL
XFILL_10_MUX2X1_180 gnd vdd FILL
XFILL_23_7 gnd vdd FILL
XFILL_62_DFFSR_12 gnd vdd FILL
XFILL_62_DFFSR_23 gnd vdd FILL
XFILL_10_MUX2X1_191 gnd vdd FILL
XFILL_22_DFFSR_210 gnd vdd FILL
XFILL_62_DFFSR_34 gnd vdd FILL
XFILL_22_DFFSR_221 gnd vdd FILL
XFILL_62_DFFSR_45 gnd vdd FILL
XFILL_3_AOI22X1_6 gnd vdd FILL
XFILL_62_DFFSR_56 gnd vdd FILL
XFILL_22_DFFSR_232 gnd vdd FILL
XFILL_16_6 gnd vdd FILL
XFILL_22_DFFSR_243 gnd vdd FILL
XFILL_15_OAI21X1_9 gnd vdd FILL
XFILL_62_DFFSR_67 gnd vdd FILL
XFILL_62_DFFSR_78 gnd vdd FILL
XFILL_22_DFFSR_254 gnd vdd FILL
XFILL_62_DFFSR_89 gnd vdd FILL
XFILL_22_DFFSR_265 gnd vdd FILL
XFILL_3_INVX1_205 gnd vdd FILL
XFILL_3_INVX1_216 gnd vdd FILL
XFILL_26_CLKBUF1_15 gnd vdd FILL
XDFFSR_6 DFFSR_6/Q DFFSR_6/CLK DFFSR_6/R vdd DFFSR_6/D gnd vdd DFFSR
XFILL_5_DFFSR_14 gnd vdd FILL
XFILL_3_INVX1_227 gnd vdd FILL
XFILL_26_CLKBUF1_26 gnd vdd FILL
XFILL_5_DFFSR_25 gnd vdd FILL
XFILL_26_DFFSR_220 gnd vdd FILL
XFILL_26_CLKBUF1_37 gnd vdd FILL
XFILL_31_DFFSR_11 gnd vdd FILL
XFILL_5_DFFSR_36 gnd vdd FILL
XFILL_7_AOI22X1_5 gnd vdd FILL
XFILL_26_DFFSR_231 gnd vdd FILL
XFILL_26_DFFSR_242 gnd vdd FILL
XFILL_5_DFFSR_47 gnd vdd FILL
XFILL_31_DFFSR_22 gnd vdd FILL
XFILL_26_DFFSR_253 gnd vdd FILL
XFILL_5_DFFSR_58 gnd vdd FILL
XFILL_31_DFFSR_33 gnd vdd FILL
XFILL_5_DFFSR_69 gnd vdd FILL
XFILL_26_DFFSR_264 gnd vdd FILL
XFILL_31_DFFSR_44 gnd vdd FILL
XFILL_9_CLKBUF1_19 gnd vdd FILL
XFILL_26_DFFSR_275 gnd vdd FILL
XFILL_31_DFFSR_55 gnd vdd FILL
XFILL_31_DFFSR_66 gnd vdd FILL
XFILL_7_INVX1_204 gnd vdd FILL
XFILL_7_INVX1_215 gnd vdd FILL
XFILL_31_DFFSR_77 gnd vdd FILL
XFILL_53_DFFSR_120 gnd vdd FILL
XFILL_7_INVX1_226 gnd vdd FILL
XFILL_53_DFFSR_131 gnd vdd FILL
XFILL_4_AOI21X1_16 gnd vdd FILL
XFILL_31_DFFSR_88 gnd vdd FILL
XFILL_31_DFFSR_99 gnd vdd FILL
XFILL_7_INVX1_90 gnd vdd FILL
XFILL_4_AOI21X1_27 gnd vdd FILL
XFILL_71_DFFSR_10 gnd vdd FILL
XFILL_71_DFFSR_21 gnd vdd FILL
XFILL_53_DFFSR_142 gnd vdd FILL
XFILL_4_AOI21X1_38 gnd vdd FILL
XFILL_7_BUFX2_10 gnd vdd FILL
XFILL_4_AOI21X1_49 gnd vdd FILL
XFILL_53_DFFSR_153 gnd vdd FILL
XFILL_71_DFFSR_32 gnd vdd FILL
XFILL_53_DFFSR_164 gnd vdd FILL
XFILL_71_DFFSR_43 gnd vdd FILL
XFILL_53_DFFSR_175 gnd vdd FILL
XFILL_14_OAI22X1_18 gnd vdd FILL
XFILL_14_OAI22X1_29 gnd vdd FILL
XFILL_71_DFFSR_54 gnd vdd FILL
XFILL_53_DFFSR_186 gnd vdd FILL
XFILL_71_DFFSR_65 gnd vdd FILL
XFILL_71_DFFSR_76 gnd vdd FILL
XFILL_53_DFFSR_197 gnd vdd FILL
XFILL_7_NOR2X1_104 gnd vdd FILL
XFILL_57_DFFSR_130 gnd vdd FILL
XFILL_71_DFFSR_87 gnd vdd FILL
XFILL_7_NOR2X1_115 gnd vdd FILL
XFILL_71_DFFSR_98 gnd vdd FILL
XFILL_7_NOR2X1_126 gnd vdd FILL
XFILL_7_NOR2X1_137 gnd vdd FILL
XFILL_57_DFFSR_141 gnd vdd FILL
XFILL_57_DFFSR_152 gnd vdd FILL
XFILL_57_DFFSR_163 gnd vdd FILL
XFILL_7_NOR2X1_148 gnd vdd FILL
XFILL_7_NOR2X1_159 gnd vdd FILL
XFILL_57_DFFSR_174 gnd vdd FILL
XNAND2X1_40 NOR2X1_45/B INVX1_138/Y gnd NOR3X1_6/C vdd NAND2X1
XFILL_0_DFFSR_101 gnd vdd FILL
XFILL_13_NAND3X1_50 gnd vdd FILL
XFILL_57_DFFSR_185 gnd vdd FILL
XNAND2X1_51 BUFX4_92/Y NOR3X1_2/Y gnd OAI21X1_3/B vdd NAND2X1
XFILL_40_DFFSR_20 gnd vdd FILL
XFILL_0_DFFSR_112 gnd vdd FILL
XFILL_13_NAND3X1_61 gnd vdd FILL
XNAND2X1_62 BUFX4_5/Y NOR2X1_30/Y gnd NOR2X1_66/B vdd NAND2X1
XFILL_40_DFFSR_31 gnd vdd FILL
XFILL_0_DFFSR_123 gnd vdd FILL
XFILL_57_DFFSR_196 gnd vdd FILL
XNAND2X1_73 NOR2X1_93/Y NOR2X1_92/Y gnd NOR3X1_35/C vdd NAND2X1
XFILL_13_NAND3X1_72 gnd vdd FILL
XFILL_11_NOR3X1_6 gnd vdd FILL
XFILL_0_DFFSR_134 gnd vdd FILL
XFILL_37_4_0 gnd vdd FILL
XFILL_13_NAND3X1_83 gnd vdd FILL
XFILL_40_DFFSR_42 gnd vdd FILL
XNAND2X1_84 INVX1_137/A INVX1_134/Y gnd OAI21X1_35/A vdd NAND2X1
XFILL_13_NAND3X1_94 gnd vdd FILL
XFILL_0_DFFSR_145 gnd vdd FILL
XFILL_40_DFFSR_53 gnd vdd FILL
XNAND2X1_95 INVX2_3/Y NOR2X1_13/B gnd NOR2X1_138/A vdd NAND2X1
XFILL_0_DFFSR_156 gnd vdd FILL
XFILL_40_DFFSR_64 gnd vdd FILL
XFILL_0_DFFSR_167 gnd vdd FILL
XFILL_40_DFFSR_75 gnd vdd FILL
XFILL_40_DFFSR_86 gnd vdd FILL
XFILL_0_DFFSR_178 gnd vdd FILL
XFILL_4_DFFSR_100 gnd vdd FILL
XFILL_0_DFFSR_189 gnd vdd FILL
XFILL_40_DFFSR_97 gnd vdd FILL
XFILL_4_DFFSR_111 gnd vdd FILL
XFILL_35_DFFSR_109 gnd vdd FILL
XFILL_80_DFFSR_30 gnd vdd FILL
XFILL_4_DFFSR_122 gnd vdd FILL
XFILL_4_DFFSR_133 gnd vdd FILL
XFILL_80_DFFSR_41 gnd vdd FILL
XFILL_4_DFFSR_144 gnd vdd FILL
XFILL_80_DFFSR_52 gnd vdd FILL
XFILL_80_DFFSR_63 gnd vdd FILL
XFILL_4_DFFSR_155 gnd vdd FILL
XFILL_80_DFFSR_74 gnd vdd FILL
XFILL_4_DFFSR_166 gnd vdd FILL
XFILL_4_DFFSR_177 gnd vdd FILL
XFILL_80_DFFSR_85 gnd vdd FILL
XFILL_80_DFFSR_96 gnd vdd FILL
XFILL_4_DFFSR_188 gnd vdd FILL
XFILL_8_DFFSR_110 gnd vdd FILL
XFILL_4_DFFSR_199 gnd vdd FILL
XFILL_7_NOR2X1_1 gnd vdd FILL
XFILL_39_DFFSR_108 gnd vdd FILL
XFILL_8_DFFSR_121 gnd vdd FILL
XFILL_8_DFFSR_132 gnd vdd FILL
XFILL_12_MUX2X1_30 gnd vdd FILL
XFILL_39_DFFSR_119 gnd vdd FILL
XFILL_8_DFFSR_143 gnd vdd FILL
XFILL_12_MUX2X1_41 gnd vdd FILL
XFILL_20_3_0 gnd vdd FILL
XFILL_8_DFFSR_154 gnd vdd FILL
XFILL_12_MUX2X1_52 gnd vdd FILL
XFILL_8_DFFSR_165 gnd vdd FILL
XFILL_12_MUX2X1_63 gnd vdd FILL
XFILL_4_OAI22X1_13 gnd vdd FILL
XFILL_12_MUX2X1_74 gnd vdd FILL
XFILL_8_DFFSR_176 gnd vdd FILL
XFILL_20_NOR3X1_4 gnd vdd FILL
XFILL_4_OAI22X1_24 gnd vdd FILL
XFILL_12_MUX2X1_85 gnd vdd FILL
XFILL_4_OAI22X1_35 gnd vdd FILL
XFILL_8_DFFSR_187 gnd vdd FILL
XFILL_0_NOR3X1_12 gnd vdd FILL
XFILL_4_OAI22X1_46 gnd vdd FILL
XFILL_0_NOR3X1_23 gnd vdd FILL
XFILL_0_NOR3X1_34 gnd vdd FILL
XFILL_12_MUX2X1_96 gnd vdd FILL
XFILL_8_DFFSR_198 gnd vdd FILL
XFILL_8_OAI21X1_15 gnd vdd FILL
XFILL_0_NOR3X1_45 gnd vdd FILL
XFILL_8_OAI21X1_26 gnd vdd FILL
XFILL_16_MUX2X1_40 gnd vdd FILL
XFILL_8_OAI21X1_37 gnd vdd FILL
XFILL_16_MUX2X1_51 gnd vdd FILL
XFILL_8_OAI21X1_48 gnd vdd FILL
XFILL_16_MUX2X1_62 gnd vdd FILL
XFILL_16_MUX2X1_73 gnd vdd FILL
XFILL_4_NOR3X1_11 gnd vdd FILL
XFILL_16_MUX2X1_84 gnd vdd FILL
XFILL_4_NOR3X1_22 gnd vdd FILL
XFILL_4_NOR3X1_33 gnd vdd FILL
XFILL_16_MUX2X1_95 gnd vdd FILL
XFILL_41_DFFSR_1 gnd vdd FILL
XFILL_4_NOR3X1_44 gnd vdd FILL
XFILL_20_DFFSR_120 gnd vdd FILL
XFILL_1_NOR2X1_204 gnd vdd FILL
XFILL_85_DFFSR_209 gnd vdd FILL
XFILL_20_DFFSR_131 gnd vdd FILL
XFILL_20_DFFSR_142 gnd vdd FILL
XFILL_7_NAND2X1_80 gnd vdd FILL
XFILL_8_NOR3X1_10 gnd vdd FILL
XFILL_20_DFFSR_153 gnd vdd FILL
XFILL_7_NAND2X1_91 gnd vdd FILL
XFILL_20_DFFSR_164 gnd vdd FILL
XFILL_20_DFFSR_175 gnd vdd FILL
XFILL_3_NOR3X1_5 gnd vdd FILL
XFILL_8_NOR3X1_21 gnd vdd FILL
XFILL_1_INVX1_104 gnd vdd FILL
XFILL_8_NOR3X1_32 gnd vdd FILL
XFILL_1_INVX1_115 gnd vdd FILL
XFILL_59_0_2 gnd vdd FILL
XFILL_20_DFFSR_186 gnd vdd FILL
XFILL_8_NOR3X1_43 gnd vdd FILL
XFILL_15_CLKBUF1_11 gnd vdd FILL
XFILL_1_INVX1_126 gnd vdd FILL
XFILL_20_DFFSR_197 gnd vdd FILL
XFILL_15_CLKBUF1_22 gnd vdd FILL
XFILL_4_BUFX2_6 gnd vdd FILL
XFILL_24_DFFSR_130 gnd vdd FILL
XFILL_15_CLKBUF1_33 gnd vdd FILL
XFILL_1_INVX1_137 gnd vdd FILL
XFILL_1_INVX1_148 gnd vdd FILL
XFILL_1_INVX1_159 gnd vdd FILL
XFILL_24_DFFSR_141 gnd vdd FILL
XFILL_24_DFFSR_152 gnd vdd FILL
XFILL_10_AOI21X1_30 gnd vdd FILL
XFILL_24_DFFSR_163 gnd vdd FILL
XFILL_24_DFFSR_174 gnd vdd FILL
XFILL_10_AOI21X1_41 gnd vdd FILL
XFILL_3_4_0 gnd vdd FILL
XFILL_5_INVX1_103 gnd vdd FILL
XFILL_24_DFFSR_185 gnd vdd FILL
XFILL_28_4_0 gnd vdd FILL
XFILL_5_INVX1_114 gnd vdd FILL
XFILL_10_AOI21X1_52 gnd vdd FILL
XFILL_5_INVX1_125 gnd vdd FILL
XFILL_10_AOI21X1_63 gnd vdd FILL
XFILL_24_DFFSR_196 gnd vdd FILL
XFILL_10_AOI21X1_74 gnd vdd FILL
XFILL_1_DFFSR_40 gnd vdd FILL
XFILL_5_INVX1_136 gnd vdd FILL
XFILL_5_INVX1_147 gnd vdd FILL
XFILL_1_DFFSR_51 gnd vdd FILL
XFILL_28_DFFSR_140 gnd vdd FILL
XFILL_1_DFFSR_62 gnd vdd FILL
XFILL_5_INVX1_158 gnd vdd FILL
XFILL_63_DFFSR_5 gnd vdd FILL
XFILL_5_INVX1_169 gnd vdd FILL
XFILL_28_DFFSR_151 gnd vdd FILL
XFILL_28_DFFSR_162 gnd vdd FILL
XFILL_1_DFFSR_73 gnd vdd FILL
XFILL_1_DFFSR_84 gnd vdd FILL
XFILL_28_DFFSR_173 gnd vdd FILL
XFILL_28_DFFSR_184 gnd vdd FILL
XFILL_1_DFFSR_95 gnd vdd FILL
XFILL_20_NOR3X1_20 gnd vdd FILL
XFILL_20_NOR3X1_31 gnd vdd FILL
XFILL_28_DFFSR_195 gnd vdd FILL
XFILL_20_NOR3X1_42 gnd vdd FILL
XFILL_70_DFFSR_220 gnd vdd FILL
XFILL_70_DFFSR_231 gnd vdd FILL
XFILL_70_DFFSR_242 gnd vdd FILL
XFILL_12_NAND3X1_102 gnd vdd FILL
XFILL_12_NAND3X1_113 gnd vdd FILL
XFILL_70_DFFSR_253 gnd vdd FILL
XFILL_12_NAND3X1_124 gnd vdd FILL
XFILL_11_3_0 gnd vdd FILL
XFILL_70_DFFSR_264 gnd vdd FILL
XFILL_70_DFFSR_275 gnd vdd FILL
XFILL_24_NOR3X1_30 gnd vdd FILL
XFILL_24_NOR3X1_41 gnd vdd FILL
XFILL_24_NOR3X1_52 gnd vdd FILL
XFILL_74_DFFSR_230 gnd vdd FILL
XFILL_3_OAI22X1_9 gnd vdd FILL
XFILL_74_DFFSR_241 gnd vdd FILL
XFILL_74_DFFSR_252 gnd vdd FILL
XFILL_28_DFFSR_8 gnd vdd FILL
XFILL_74_DFFSR_263 gnd vdd FILL
XFILL_74_DFFSR_274 gnd vdd FILL
XFILL_28_NOR3X1_40 gnd vdd FILL
XFILL_85_DFFSR_9 gnd vdd FILL
XFILL_28_NOR3X1_51 gnd vdd FILL
XFILL_13_MUX2X1_102 gnd vdd FILL
XFILL_13_MUX2X1_113 gnd vdd FILL
XFILL_13_MUX2X1_124 gnd vdd FILL
XFILL_7_OAI22X1_8 gnd vdd FILL
XFILL_13_MUX2X1_135 gnd vdd FILL
XFILL_3_NAND3X1_107 gnd vdd FILL
XFILL_78_DFFSR_240 gnd vdd FILL
XFILL_13_MUX2X1_146 gnd vdd FILL
XFILL_3_NAND3X1_118 gnd vdd FILL
XFILL_78_DFFSR_251 gnd vdd FILL
XFILL_3_NAND3X1_129 gnd vdd FILL
XFILL_78_DFFSR_262 gnd vdd FILL
XFILL_13_MUX2X1_157 gnd vdd FILL
XFILL_33_CLKBUF1_3 gnd vdd FILL
XFILL_13_MUX2X1_168 gnd vdd FILL
XFILL_78_DFFSR_273 gnd vdd FILL
XFILL_0_AOI21X1_80 gnd vdd FILL
XFILL_13_MUX2X1_179 gnd vdd FILL
XFILL_52_DFFSR_209 gnd vdd FILL
XFILL_14_OAI21X1_40 gnd vdd FILL
XFILL_2_INVX1_4 gnd vdd FILL
XFILL_3_NOR2X1_190 gnd vdd FILL
XFILL_56_DFFSR_208 gnd vdd FILL
XFILL_56_DFFSR_219 gnd vdd FILL
XFILL_19_4_0 gnd vdd FILL
XFILL_62_7_1 gnd vdd FILL
XFILL_83_DFFSR_108 gnd vdd FILL
XFILL_83_DFFSR_119 gnd vdd FILL
XFILL_61_2_0 gnd vdd FILL
XFILL_21_4 gnd vdd FILL
XFILL_20_MUX2X1_170 gnd vdd FILL
XFILL_20_MUX2X1_181 gnd vdd FILL
XFILL_87_DFFSR_107 gnd vdd FILL
XFILL_14_3 gnd vdd FILL
XFILL_20_MUX2X1_192 gnd vdd FILL
XFILL_87_DFFSR_118 gnd vdd FILL
XFILL_3_MUX2X1_130 gnd vdd FILL
XFILL_14_BUFX4_12 gnd vdd FILL
XFILL_3_MUX2X1_141 gnd vdd FILL
XFILL_87_DFFSR_129 gnd vdd FILL
XFILL_3_MUX2X1_152 gnd vdd FILL
XFILL_14_BUFX4_23 gnd vdd FILL
XFILL_3_MUX2X1_163 gnd vdd FILL
XFILL_14_BUFX4_34 gnd vdd FILL
XFILL_14_BUFX4_45 gnd vdd FILL
XFILL_3_MUX2X1_174 gnd vdd FILL
XDFFSR_202 INVX1_94/A DFFSR_45/CLK DFFSR_57/R vdd MUX2X1_81/Y gnd vdd DFFSR
XFILL_3_MUX2X1_185 gnd vdd FILL
XFILL_14_BUFX4_56 gnd vdd FILL
XDFFSR_213 INVX1_88/A DFFSR_57/CLK DFFSR_57/R vdd MUX2X1_75/Y gnd vdd DFFSR
XFILL_14_BUFX4_67 gnd vdd FILL
XFILL_14_BUFX4_78 gnd vdd FILL
XDFFSR_224 INVX1_73/A CLKBUF1_26/Y DFFSR_25/R vdd MUX2X1_60/Y gnd vdd DFFSR
XDFFSR_235 INVX1_66/A DFFSR_4/CLK DFFSR_23/R vdd MUX2X1_53/Y gnd vdd DFFSR
XFILL_14_BUFX4_89 gnd vdd FILL
XDFFSR_246 INVX1_51/A DFFSR_39/CLK BUFX4_50/Y vdd MUX2X1_38/Y gnd vdd DFFSR
XDFFSR_257 NOR2X1_19/A DFFSR_5/CLK DFFSR_5/R vdd DFFSR_257/D gnd vdd DFFSR
XDFFSR_268 INVX1_37/A DFFSR_5/CLK DFFSR_5/R vdd MUX2X1_23/Y gnd vdd DFFSR
XFILL_41_DFFSR_230 gnd vdd FILL
XFILL_41_DFFSR_241 gnd vdd FILL
XFILL_41_DFFSR_252 gnd vdd FILL
XFILL_41_DFFSR_263 gnd vdd FILL
XFILL_41_DFFSR_274 gnd vdd FILL
XFILL_8_NAND3X1_9 gnd vdd FILL
XFILL_45_DFFSR_240 gnd vdd FILL
XFILL_45_DFFSR_251 gnd vdd FILL
XFILL_45_DFFSR_262 gnd vdd FILL
XFILL_45_DFFSR_273 gnd vdd FILL
XFILL_72_DFFSR_140 gnd vdd FILL
XFILL_9_AND2X2_5 gnd vdd FILL
XFILL_72_DFFSR_151 gnd vdd FILL
XFILL_49_DFFSR_250 gnd vdd FILL
XFILL_72_DFFSR_162 gnd vdd FILL
XFILL_49_DFFSR_261 gnd vdd FILL
XFILL_72_DFFSR_173 gnd vdd FILL
XFILL_72_DFFSR_184 gnd vdd FILL
XFILL_49_DFFSR_272 gnd vdd FILL
XFILL_72_DFFSR_195 gnd vdd FILL
XFILL_23_DFFSR_208 gnd vdd FILL
XFILL_6_NAND3X1_11 gnd vdd FILL
XFILL_6_NAND3X1_22 gnd vdd FILL
XFILL_23_DFFSR_219 gnd vdd FILL
XFILL_6_NAND3X1_33 gnd vdd FILL
XFILL_53_7_1 gnd vdd FILL
XFILL_76_DFFSR_150 gnd vdd FILL
XFILL_6_NAND3X1_44 gnd vdd FILL
XFILL_76_DFFSR_161 gnd vdd FILL
XFILL_6_NAND3X1_55 gnd vdd FILL
XFILL_6_NAND3X1_66 gnd vdd FILL
XFILL_76_DFFSR_172 gnd vdd FILL
XFILL_45_DFFSR_2 gnd vdd FILL
XFILL_6_NAND3X1_77 gnd vdd FILL
XFILL_6_BUFX4_11 gnd vdd FILL
XFILL_52_2_0 gnd vdd FILL
XFILL_76_DFFSR_183 gnd vdd FILL
XFILL_6_BUFX4_22 gnd vdd FILL
XFILL_76_DFFSR_194 gnd vdd FILL
XFILL_50_DFFSR_108 gnd vdd FILL
XFILL_6_BUFX4_33 gnd vdd FILL
XFILL_6_NAND3X1_88 gnd vdd FILL
XFILL_27_DFFSR_207 gnd vdd FILL
XFILL_6_NAND3X1_99 gnd vdd FILL
XFILL_50_DFFSR_119 gnd vdd FILL
XFILL_6_BUFX4_44 gnd vdd FILL
XFILL_27_DFFSR_218 gnd vdd FILL
XFILL_27_DFFSR_229 gnd vdd FILL
XFILL_6_BUFX4_55 gnd vdd FILL
XFILL_6_BUFX4_66 gnd vdd FILL
XFILL_6_BUFX4_77 gnd vdd FILL
XFILL_6_BUFX4_88 gnd vdd FILL
XFILL_6_BUFX4_99 gnd vdd FILL
XFILL_54_DFFSR_107 gnd vdd FILL
XFILL_8_BUFX2_7 gnd vdd FILL
XFILL_54_DFFSR_118 gnd vdd FILL
XFILL_54_DFFSR_129 gnd vdd FILL
XFILL_81_DFFSR_19 gnd vdd FILL
XFILL_13_AOI21X1_18 gnd vdd FILL
XFILL_13_AOI21X1_29 gnd vdd FILL
XFILL_10_DFFSR_19 gnd vdd FILL
XFILL_58_DFFSR_106 gnd vdd FILL
XFILL_58_DFFSR_117 gnd vdd FILL
XFILL_58_DFFSR_128 gnd vdd FILL
XFILL_58_DFFSR_139 gnd vdd FILL
XFILL_67_DFFSR_6 gnd vdd FILL
XFILL_50_DFFSR_18 gnd vdd FILL
XFILL_50_DFFSR_29 gnd vdd FILL
XFILL_7_0_2 gnd vdd FILL
XFILL_12_DFFSR_240 gnd vdd FILL
XFILL_12_DFFSR_251 gnd vdd FILL
XFILL_12_DFFSR_262 gnd vdd FILL
XFILL_5_DFFSR_109 gnd vdd FILL
XFILL_12_DFFSR_273 gnd vdd FILL
XFILL_25_CLKBUF1_12 gnd vdd FILL
XFILL_25_CLKBUF1_23 gnd vdd FILL
XFILL_25_CLKBUF1_34 gnd vdd FILL
XFILL_0_AOI21X1_5 gnd vdd FILL
XFILL_10_BUFX4_60 gnd vdd FILL
XFILL_16_DFFSR_250 gnd vdd FILL
XFILL_10_BUFX4_71 gnd vdd FILL
XFILL_7_BUFX4_1 gnd vdd FILL
XFILL_16_DFFSR_261 gnd vdd FILL
XFILL_10_BUFX4_82 gnd vdd FILL
XFILL_9_DFFSR_108 gnd vdd FILL
XFILL_8_CLKBUF1_16 gnd vdd FILL
XFILL_16_DFFSR_272 gnd vdd FILL
XFILL_10_BUFX4_93 gnd vdd FILL
XFILL_9_DFFSR_119 gnd vdd FILL
XFILL_13_MUX2X1_17 gnd vdd FILL
XFILL_8_CLKBUF1_27 gnd vdd FILL
XFILL_8_CLKBUF1_38 gnd vdd FILL
XFILL_44_7_1 gnd vdd FILL
XFILL_13_MUX2X1_28 gnd vdd FILL
XFILL_3_AOI21X1_13 gnd vdd FILL
XFILL_13_MUX2X1_39 gnd vdd FILL
XFILL_43_2_0 gnd vdd FILL
XFILL_3_AOI21X1_24 gnd vdd FILL
XFILL_4_AOI21X1_4 gnd vdd FILL
XFILL_3_AOI21X1_35 gnd vdd FILL
XFILL_3_AOI21X1_46 gnd vdd FILL
XFILL_43_DFFSR_150 gnd vdd FILL
XFILL_43_DFFSR_161 gnd vdd FILL
XFILL_3_AOI21X1_57 gnd vdd FILL
XOAI21X1_16 INVX1_193/Y OAI21X1_6/B OAI21X1_16/C gnd NOR2X1_78/B vdd OAI21X1
XFILL_43_DFFSR_172 gnd vdd FILL
XFILL_13_OAI22X1_15 gnd vdd FILL
XFILL_3_AOI21X1_68 gnd vdd FILL
XFILL_43_DFFSR_183 gnd vdd FILL
XFILL_13_OAI22X1_26 gnd vdd FILL
XOAI21X1_27 INVX1_169/Y OAI21X1_2/B OAI21X1_27/C gnd OAI21X1_27/Y vdd OAI21X1
XFILL_17_MUX2X1_16 gnd vdd FILL
XFILL_3_AOI21X1_79 gnd vdd FILL
XFILL_13_OAI22X1_37 gnd vdd FILL
XFILL_43_DFFSR_194 gnd vdd FILL
XOAI21X1_38 BUFX2_9/A AND2X2_8/B OAI21X1_38/C gnd OAI21X1_1/C vdd OAI21X1
XFILL_17_MUX2X1_27 gnd vdd FILL
XOAI21X1_49 NOR3X1_2/Y AND2X2_1/Y BUFX4_60/Y gnd OAI21X1_49/Y vdd OAI21X1
XFILL_6_NOR2X1_101 gnd vdd FILL
XFILL_17_MUX2X1_38 gnd vdd FILL
XFILL_13_OAI22X1_48 gnd vdd FILL
XFILL_8_AOI21X1_3 gnd vdd FILL
XFILL_6_NOR2X1_112 gnd vdd FILL
XFILL_6_NOR2X1_123 gnd vdd FILL
XFILL_17_MUX2X1_49 gnd vdd FILL
XFILL_6_NOR2X1_134 gnd vdd FILL
XFILL_6_NOR2X1_145 gnd vdd FILL
XFILL_13_NAND3X1_103 gnd vdd FILL
XFILL_2_DFFSR_18 gnd vdd FILL
XFILL_47_DFFSR_160 gnd vdd FILL
XFILL_2_DFFSR_29 gnd vdd FILL
XFILL_13_NAND3X1_114 gnd vdd FILL
XFILL_6_NOR2X1_156 gnd vdd FILL
XFILL_47_DFFSR_171 gnd vdd FILL
XFILL_6_INVX1_5 gnd vdd FILL
XFILL_13_NAND3X1_125 gnd vdd FILL
XFILL_6_NOR2X1_167 gnd vdd FILL
XFILL_47_DFFSR_182 gnd vdd FILL
XFILL_6_NOR2X1_178 gnd vdd FILL
XFILL_47_DFFSR_193 gnd vdd FILL
XFILL_21_DFFSR_107 gnd vdd FILL
XFILL_6_NOR2X1_189 gnd vdd FILL
XFILL_21_DFFSR_118 gnd vdd FILL
XFILL_4_INVX1_50 gnd vdd FILL
XFILL_12_NAND3X1_80 gnd vdd FILL
XFILL_21_DFFSR_129 gnd vdd FILL
XFILL_12_NAND3X1_91 gnd vdd FILL
XFILL_4_INVX1_61 gnd vdd FILL
XFILL_10_NOR2X1_206 gnd vdd FILL
XFILL_4_INVX1_72 gnd vdd FILL
XFILL_4_INVX1_83 gnd vdd FILL
XFILL_9_NOR3X1_19 gnd vdd FILL
XFILL_4_INVX1_94 gnd vdd FILL
XFILL_25_DFFSR_106 gnd vdd FILL
XFILL_25_DFFSR_117 gnd vdd FILL
XFILL_11_MUX2X1_4 gnd vdd FILL
XFILL_23_MUX2X1_103 gnd vdd FILL
XFILL_25_DFFSR_128 gnd vdd FILL
XFILL_23_MUX2X1_114 gnd vdd FILL
XFILL_23_MUX2X1_125 gnd vdd FILL
XFILL_25_DFFSR_139 gnd vdd FILL
XFILL_23_MUX2X1_136 gnd vdd FILL
XFILL_4_NAND3X1_108 gnd vdd FILL
XFILL_4_NAND3X1_119 gnd vdd FILL
XFILL_23_MUX2X1_147 gnd vdd FILL
XFILL_23_MUX2X1_158 gnd vdd FILL
XFILL_23_MUX2X1_169 gnd vdd FILL
XFILL_7_INVX4_1 gnd vdd FILL
XFILL_6_MUX2X1_107 gnd vdd FILL
XFILL_29_DFFSR_105 gnd vdd FILL
XFILL_6_MUX2X1_118 gnd vdd FILL
XFILL_29_DFFSR_116 gnd vdd FILL
XFILL_6_MUX2X1_129 gnd vdd FILL
XFILL_29_DFFSR_127 gnd vdd FILL
XFILL_19_DFFSR_30 gnd vdd FILL
XFILL_29_DFFSR_138 gnd vdd FILL
XFILL_2_BUFX4_70 gnd vdd FILL
XFILL_19_DFFSR_41 gnd vdd FILL
XFILL_2_BUFX4_81 gnd vdd FILL
XFILL_29_DFFSR_149 gnd vdd FILL
XFILL_2_BUFX4_92 gnd vdd FILL
XFILL_3_OAI22X1_10 gnd vdd FILL
XFILL_19_DFFSR_52 gnd vdd FILL
XFILL_19_DFFSR_63 gnd vdd FILL
XFILL_3_OAI22X1_21 gnd vdd FILL
XFILL_19_DFFSR_74 gnd vdd FILL
XFILL_3_OAI22X1_32 gnd vdd FILL
XFILL_3_OAI22X1_43 gnd vdd FILL
XFILL_19_DFFSR_85 gnd vdd FILL
XFILL_21_NOR3X1_18 gnd vdd FILL
XFILL_19_DFFSR_96 gnd vdd FILL
XFILL_7_OAI21X1_12 gnd vdd FILL
XFILL_21_NOR3X1_29 gnd vdd FILL
XFILL_7_OAI21X1_23 gnd vdd FILL
XFILL_7_OAI21X1_34 gnd vdd FILL
XFILL_71_DFFSR_207 gnd vdd FILL
XFILL_59_DFFSR_40 gnd vdd FILL
XFILL_59_DFFSR_51 gnd vdd FILL
XFILL_71_DFFSR_218 gnd vdd FILL
XFILL_7_OAI21X1_45 gnd vdd FILL
XFILL_71_DFFSR_229 gnd vdd FILL
XFILL_20_MUX2X1_2 gnd vdd FILL
XFILL_35_7_1 gnd vdd FILL
XFILL_59_DFFSR_62 gnd vdd FILL
XFILL_59_DFFSR_73 gnd vdd FILL
XFILL_59_DFFSR_84 gnd vdd FILL
XFILL_59_DFFSR_95 gnd vdd FILL
XFILL_25_NOR3X1_17 gnd vdd FILL
XFILL_34_2_0 gnd vdd FILL
XFILL_25_NOR3X1_28 gnd vdd FILL
XFILL_25_NOR3X1_39 gnd vdd FILL
XFILL_75_DFFSR_206 gnd vdd FILL
XFILL_0_NOR2X1_201 gnd vdd FILL
XFILL_4_NOR2X1_5 gnd vdd FILL
XFILL_75_DFFSR_217 gnd vdd FILL
XFILL_75_DFFSR_228 gnd vdd FILL
XFILL_10_DFFSR_150 gnd vdd FILL
XFILL_75_DFFSR_239 gnd vdd FILL
XFILL_10_DFFSR_161 gnd vdd FILL
XFILL_29_NOR3X1_16 gnd vdd FILL
XFILL_10_DFFSR_172 gnd vdd FILL
XFILL_10_DFFSR_183 gnd vdd FILL
XFILL_28_DFFSR_50 gnd vdd FILL
XFILL_29_NOR3X1_27 gnd vdd FILL
XFILL_28_DFFSR_61 gnd vdd FILL
XFILL_29_NOR3X1_38 gnd vdd FILL
XFILL_10_DFFSR_194 gnd vdd FILL
XFILL_29_NOR3X1_49 gnd vdd FILL
XFILL_79_DFFSR_205 gnd vdd FILL
XFILL_28_DFFSR_72 gnd vdd FILL
XFILL_28_DFFSR_83 gnd vdd FILL
XFILL_14_CLKBUF1_30 gnd vdd FILL
XFILL_14_CLKBUF1_41 gnd vdd FILL
XFILL_79_DFFSR_216 gnd vdd FILL
XFILL_28_DFFSR_94 gnd vdd FILL
XFILL_79_DFFSR_227 gnd vdd FILL
XFILL_79_DFFSR_238 gnd vdd FILL
XFILL_14_DFFSR_160 gnd vdd FILL
XFILL_79_DFFSR_249 gnd vdd FILL
XFILL_3_CLKBUF1_3 gnd vdd FILL
XFILL_3_MUX2X1_3 gnd vdd FILL
XFILL_14_DFFSR_171 gnd vdd FILL
XFILL_14_DFFSR_182 gnd vdd FILL
XFILL_14_DFFSR_193 gnd vdd FILL
XFILL_68_DFFSR_60 gnd vdd FILL
XFILL_68_DFFSR_71 gnd vdd FILL
XFILL_68_DFFSR_82 gnd vdd FILL
XFILL_11_DFFSR_5 gnd vdd FILL
XFILL_68_DFFSR_93 gnd vdd FILL
XFILL_49_DFFSR_3 gnd vdd FILL
XFILL_18_DFFSR_170 gnd vdd FILL
XFILL_7_CLKBUF1_2 gnd vdd FILL
XFILL_18_DFFSR_181 gnd vdd FILL
XFILL_18_DFFSR_192 gnd vdd FILL
XFILL_0_NOR3X1_9 gnd vdd FILL
XFILL_10_NOR3X1_50 gnd vdd FILL
XFILL_37_DFFSR_70 gnd vdd FILL
XFILL_37_DFFSR_81 gnd vdd FILL
XFILL_60_DFFSR_250 gnd vdd FILL
XFILL_37_DFFSR_92 gnd vdd FILL
XFILL_60_DFFSR_261 gnd vdd FILL
XFILL_60_DFFSR_272 gnd vdd FILL
XFILL_77_DFFSR_80 gnd vdd FILL
XFILL_77_DFFSR_91 gnd vdd FILL
XFILL_64_DFFSR_260 gnd vdd FILL
XFILL_33_DFFSR_9 gnd vdd FILL
XFILL_64_DFFSR_271 gnd vdd FILL
XFILL_1_7_1 gnd vdd FILL
XFILL_26_7_1 gnd vdd FILL
XFILL_12_MUX2X1_110 gnd vdd FILL
XFILL_12_MUX2X1_121 gnd vdd FILL
XFILL_25_2_0 gnd vdd FILL
XFILL_0_OAI21X1_8 gnd vdd FILL
XFILL_0_2_0 gnd vdd FILL
XFILL_12_MUX2X1_132 gnd vdd FILL
XFILL_12_MUX2X1_143 gnd vdd FILL
XFILL_12_MUX2X1_154 gnd vdd FILL
XFILL_12_MUX2X1_165 gnd vdd FILL
XFILL_68_DFFSR_270 gnd vdd FILL
XFILL_12_MUX2X1_176 gnd vdd FILL
XFILL_12_MUX2X1_187 gnd vdd FILL
XFILL_46_DFFSR_90 gnd vdd FILL
XFILL_1_NOR2X1_10 gnd vdd FILL
XFILL_42_DFFSR_206 gnd vdd FILL
XFILL_1_NOR2X1_21 gnd vdd FILL
XFILL_42_DFFSR_217 gnd vdd FILL
XFILL_1_NOR2X1_32 gnd vdd FILL
XFILL_1_NOR2X1_43 gnd vdd FILL
XFILL_4_OAI21X1_7 gnd vdd FILL
XFILL_42_DFFSR_228 gnd vdd FILL
XFILL_42_DFFSR_239 gnd vdd FILL
XFILL_1_NOR2X1_54 gnd vdd FILL
XFILL_1_NOR2X1_65 gnd vdd FILL
XFILL_1_NOR2X1_76 gnd vdd FILL
XFILL_1_NOR2X1_87 gnd vdd FILL
XFILL_46_DFFSR_205 gnd vdd FILL
XFILL_1_NOR2X1_98 gnd vdd FILL
XFILL_5_NOR2X1_20 gnd vdd FILL
XFILL_8_OAI21X1_6 gnd vdd FILL
XFILL_5_NOR2X1_31 gnd vdd FILL
XFILL_46_DFFSR_216 gnd vdd FILL
XFILL_5_NOR2X1_42 gnd vdd FILL
XFILL_46_DFFSR_227 gnd vdd FILL
XFILL_46_DFFSR_238 gnd vdd FILL
XFILL_5_NOR2X1_53 gnd vdd FILL
XFILL_46_DFFSR_249 gnd vdd FILL
XFILL_5_NOR2X1_64 gnd vdd FILL
XFILL_5_NOR2X1_75 gnd vdd FILL
XFILL_5_NOR2X1_86 gnd vdd FILL
XFILL_5_NOR2X1_97 gnd vdd FILL
XFILL_73_DFFSR_105 gnd vdd FILL
XFILL_73_DFFSR_116 gnd vdd FILL
XFILL_9_NOR2X1_30 gnd vdd FILL
XFILL_73_DFFSR_127 gnd vdd FILL
XFILL_73_DFFSR_138 gnd vdd FILL
XFILL_9_NOR2X1_41 gnd vdd FILL
XFILL_9_NOR2X1_52 gnd vdd FILL
XFILL_13_OAI22X1_3 gnd vdd FILL
XFILL_73_DFFSR_149 gnd vdd FILL
XFILL_9_NOR2X1_63 gnd vdd FILL
XFILL_9_NOR2X1_74 gnd vdd FILL
XFILL_9_NOR2X1_85 gnd vdd FILL
XFILL_8_3_0 gnd vdd FILL
XFILL_9_NOR2X1_96 gnd vdd FILL
XFILL_77_DFFSR_104 gnd vdd FILL
XFILL_6_9 gnd vdd FILL
XFILL_77_DFFSR_115 gnd vdd FILL
XFILL_77_DFFSR_126 gnd vdd FILL
XFILL_77_DFFSR_137 gnd vdd FILL
XFILL_17_OAI22X1_2 gnd vdd FILL
XFILL_2_MUX2X1_160 gnd vdd FILL
XFILL_15_NAND3X1_13 gnd vdd FILL
XFILL_77_DFFSR_148 gnd vdd FILL
XFILL_2_MUX2X1_171 gnd vdd FILL
XFILL_77_DFFSR_159 gnd vdd FILL
XFILL_15_NAND3X1_24 gnd vdd FILL
XFILL_2_MUX2X1_182 gnd vdd FILL
XFILL_15_NAND3X1_35 gnd vdd FILL
XFILL_15_NAND3X1_46 gnd vdd FILL
XFILL_2_MUX2X1_193 gnd vdd FILL
XFILL_15_NAND3X1_57 gnd vdd FILL
XFILL_15_NAND3X1_68 gnd vdd FILL
XFILL_35_CLKBUF1_13 gnd vdd FILL
XFILL_35_CLKBUF1_24 gnd vdd FILL
XFILL_15_NAND3X1_79 gnd vdd FILL
XFILL_35_CLKBUF1_35 gnd vdd FILL
XFILL_17_7_1 gnd vdd FILL
XFILL_31_DFFSR_260 gnd vdd FILL
XFILL_31_DFFSR_271 gnd vdd FILL
XFILL_16_2_0 gnd vdd FILL
XFILL_1_NAND2X1_9 gnd vdd FILL
XFILL_11_BUFX4_16 gnd vdd FILL
XFILL_11_BUFX4_27 gnd vdd FILL
XFILL_35_DFFSR_270 gnd vdd FILL
XFILL_11_BUFX4_38 gnd vdd FILL
XFILL_11_BUFX4_49 gnd vdd FILL
XFILL_5_NAND2X1_8 gnd vdd FILL
XFILL_1_MUX2X1_50 gnd vdd FILL
XFILL_1_MUX2X1_61 gnd vdd FILL
XFILL_1_MUX2X1_72 gnd vdd FILL
XFILL_1_MUX2X1_83 gnd vdd FILL
XFILL_14_NAND3X1_104 gnd vdd FILL
XFILL_1_MUX2X1_94 gnd vdd FILL
XFILL_62_DFFSR_170 gnd vdd FILL
XFILL_14_NAND3X1_115 gnd vdd FILL
XDFFSR_19 DFFSR_19/Q CLKBUF1_1/Y DFFSR_93/R vdd DFFSR_19/D gnd vdd DFFSR
XFILL_14_NAND3X1_126 gnd vdd FILL
XFILL_62_DFFSR_181 gnd vdd FILL
XFILL_62_DFFSR_192 gnd vdd FILL
XFILL_9_NAND2X1_7 gnd vdd FILL
XFILL_13_DFFSR_205 gnd vdd FILL
XFILL_10_NAND3X1_5 gnd vdd FILL
XFILL_13_DFFSR_216 gnd vdd FILL
XFILL_13_DFFSR_227 gnd vdd FILL
XFILL_5_NAND3X1_30 gnd vdd FILL
XFILL_5_MUX2X1_60 gnd vdd FILL
XFILL_5_MUX2X1_71 gnd vdd FILL
XFILL_13_DFFSR_238 gnd vdd FILL
XFILL_13_DFFSR_249 gnd vdd FILL
XFILL_5_MUX2X1_82 gnd vdd FILL
XFILL_5_NAND3X1_41 gnd vdd FILL
XFILL_50_DFFSR_3 gnd vdd FILL
XFILL_5_MUX2X1_93 gnd vdd FILL
XFILL_9_NAND2X1_10 gnd vdd FILL
XFILL_5_NAND3X1_52 gnd vdd FILL
XFILL_5_NAND3X1_63 gnd vdd FILL
XFILL_66_DFFSR_180 gnd vdd FILL
XFILL_5_NAND3X1_74 gnd vdd FILL
XFILL_9_NAND2X1_21 gnd vdd FILL
XFILL_5_NAND3X1_85 gnd vdd FILL
XFILL_9_NAND2X1_32 gnd vdd FILL
XFILL_66_DFFSR_191 gnd vdd FILL
XFILL_40_DFFSR_105 gnd vdd FILL
XFILL_17_DFFSR_204 gnd vdd FILL
XFILL_9_NAND2X1_43 gnd vdd FILL
XFILL_5_NAND3X1_96 gnd vdd FILL
XFILL_40_DFFSR_116 gnd vdd FILL
XFILL_14_NAND3X1_4 gnd vdd FILL
XFILL_9_NAND2X1_54 gnd vdd FILL
XFILL_17_DFFSR_215 gnd vdd FILL
XFILL_9_NAND2X1_65 gnd vdd FILL
XFILL_40_DFFSR_127 gnd vdd FILL
XFILL_17_DFFSR_226 gnd vdd FILL
XFILL_40_DFFSR_138 gnd vdd FILL
XFILL_17_DFFSR_237 gnd vdd FILL
XFILL_9_MUX2X1_70 gnd vdd FILL
XFILL_5_INVX1_17 gnd vdd FILL
XFILL_9_NAND2X1_76 gnd vdd FILL
XFILL_9_MUX2X1_81 gnd vdd FILL
XFILL_40_DFFSR_149 gnd vdd FILL
XFILL_17_DFFSR_248 gnd vdd FILL
XFILL_9_NAND2X1_87 gnd vdd FILL
XFILL_5_INVX1_28 gnd vdd FILL
XFILL_22_14 gnd vdd FILL
XFILL_9_MUX2X1_92 gnd vdd FILL
XFILL_5_INVX1_39 gnd vdd FILL
XFILL_17_DFFSR_259 gnd vdd FILL
XFILL_5_NAND3X1_109 gnd vdd FILL
XCLKBUF1_17 BUFX4_73/Y gnd DFFSR_97/CLK vdd CLKBUF1
XCLKBUF1_28 BUFX4_4/Y gnd DFFSR_5/CLK vdd CLKBUF1
XCLKBUF1_39 BUFX4_9/Y gnd DFFSR_57/CLK vdd CLKBUF1
XFILL_44_DFFSR_104 gnd vdd FILL
XFILL_67_1 gnd vdd FILL
XFILL_17_CLKBUF1_18 gnd vdd FILL
XFILL_44_DFFSR_115 gnd vdd FILL
XFILL_17_CLKBUF1_29 gnd vdd FILL
XFILL_44_DFFSR_126 gnd vdd FILL
XFILL_44_DFFSR_137 gnd vdd FILL
XFILL_66_1_0 gnd vdd FILL
XFILL_44_DFFSR_148 gnd vdd FILL
XBUFX4_60 BUFX4_60/A gnd BUFX4_60/Y vdd BUFX4
XFILL_12_AOI21X1_15 gnd vdd FILL
XBUFX4_71 INVX8_2/Y gnd BUFX4_71/Y vdd BUFX4
XFILL_12_AOI21X1_26 gnd vdd FILL
XFILL_44_DFFSR_159 gnd vdd FILL
XFILL_12_AOI21X1_37 gnd vdd FILL
XBUFX4_82 INVX8_4/Y gnd MUX2X1_4/B vdd BUFX4
XBUFX4_93 INVX8_3/Y gnd BUFX4_93/Y vdd BUFX4
XFILL_2_DFFSR_8 gnd vdd FILL
XFILL_12_AOI21X1_48 gnd vdd FILL
XFILL_12_AOI21X1_59 gnd vdd FILL
XFILL_48_DFFSR_103 gnd vdd FILL
XFILL_15_DFFSR_6 gnd vdd FILL
XFILL_48_DFFSR_114 gnd vdd FILL
XFILL_3_BUFX4_15 gnd vdd FILL
XFILL_48_DFFSR_125 gnd vdd FILL
XFILL_48_DFFSR_136 gnd vdd FILL
XFILL_3_BUFX4_26 gnd vdd FILL
XFILL_72_DFFSR_7 gnd vdd FILL
XFILL_3_BUFX4_37 gnd vdd FILL
XFILL_48_DFFSR_147 gnd vdd FILL
XFILL_48_DFFSR_158 gnd vdd FILL
XFILL_3_BUFX4_48 gnd vdd FILL
XFILL_21_MUX2X1_80 gnd vdd FILL
XFILL_3_BUFX4_59 gnd vdd FILL
XFILL_48_DFFSR_169 gnd vdd FILL
XFILL_21_MUX2X1_91 gnd vdd FILL
XFILL_50_5_1 gnd vdd FILL
XFILL_14_AOI22X1_9 gnd vdd FILL
XFILL_24_CLKBUF1_20 gnd vdd FILL
XFILL_24_CLKBUF1_31 gnd vdd FILL
XFILL_24_CLKBUF1_42 gnd vdd FILL
XFILL_18_AOI22X1_8 gnd vdd FILL
XFILL_0_NAND3X1_105 gnd vdd FILL
XFILL_0_NAND3X1_116 gnd vdd FILL
XFILL_63_10 gnd vdd FILL
XFILL_0_NAND3X1_127 gnd vdd FILL
XFILL_7_CLKBUF1_13 gnd vdd FILL
XFILL_7_CLKBUF1_24 gnd vdd FILL
XFILL_10_AND2X2_3 gnd vdd FILL
XFILL_29_DFFSR_17 gnd vdd FILL
XFILL_7_CLKBUF1_35 gnd vdd FILL
XFILL_2_AOI21X1_10 gnd vdd FILL
XFILL_29_DFFSR_28 gnd vdd FILL
XFILL_15_MUX2X1_109 gnd vdd FILL
XOR2X2_1 OR2X2_1/A OR2X2_1/B gnd OR2X2_1/Y vdd OR2X2
XFILL_29_DFFSR_39 gnd vdd FILL
XFILL_2_AOI21X1_21 gnd vdd FILL
XFILL_2_AOI21X1_32 gnd vdd FILL
XFILL_2_AOI21X1_43 gnd vdd FILL
XFILL_2_AOI21X1_54 gnd vdd FILL
XFILL_12_OAI22X1_12 gnd vdd FILL
XFILL_33_DFFSR_180 gnd vdd FILL
XFILL_12_OAI22X1_23 gnd vdd FILL
XFILL_2_AOI21X1_65 gnd vdd FILL
XFILL_12_OAI22X1_34 gnd vdd FILL
XFILL_2_AOI21X1_76 gnd vdd FILL
XFILL_33_DFFSR_191 gnd vdd FILL
XFILL_69_DFFSR_16 gnd vdd FILL
XFILL_12_OAI22X1_45 gnd vdd FILL
XFILL_69_DFFSR_27 gnd vdd FILL
XFILL_69_DFFSR_38 gnd vdd FILL
XFILL_69_DFFSR_49 gnd vdd FILL
XFILL_5_NOR2X1_120 gnd vdd FILL
XFILL_5_NOR2X1_131 gnd vdd FILL
XFILL_5_NOR2X1_142 gnd vdd FILL
XFILL_58_6_1 gnd vdd FILL
XFILL_5_NOR2X1_153 gnd vdd FILL
XFILL_5_NOR2X1_164 gnd vdd FILL
XFILL_57_1_0 gnd vdd FILL
XFILL_37_DFFSR_190 gnd vdd FILL
XFILL_5_NOR2X1_175 gnd vdd FILL
XFILL_11_DFFSR_104 gnd vdd FILL
XFILL_5_NOR2X1_186 gnd vdd FILL
XFILL_5_NOR2X1_197 gnd vdd FILL
XFILL_11_DFFSR_115 gnd vdd FILL
XFILL_11_DFFSR_126 gnd vdd FILL
XFILL_11_DFFSR_137 gnd vdd FILL
XFILL_38_DFFSR_15 gnd vdd FILL
XFILL_11_DFFSR_148 gnd vdd FILL
XFILL_38_DFFSR_26 gnd vdd FILL
XFILL_11_DFFSR_159 gnd vdd FILL
XFILL_38_DFFSR_37 gnd vdd FILL
XFILL_38_DFFSR_48 gnd vdd FILL
XFILL_38_DFFSR_59 gnd vdd FILL
XFILL_15_DFFSR_103 gnd vdd FILL
XFILL_15_DFFSR_114 gnd vdd FILL
XFILL_22_MUX2X1_100 gnd vdd FILL
XFILL_15_DFFSR_125 gnd vdd FILL
XFILL_15_DFFSR_136 gnd vdd FILL
XFILL_22_MUX2X1_111 gnd vdd FILL
XFILL_22_MUX2X1_122 gnd vdd FILL
XFILL_78_DFFSR_14 gnd vdd FILL
XFILL_78_DFFSR_25 gnd vdd FILL
XFILL_15_DFFSR_147 gnd vdd FILL
XFILL_22_MUX2X1_133 gnd vdd FILL
XFILL_15_DFFSR_158 gnd vdd FILL
XFILL_22_MUX2X1_144 gnd vdd FILL
XFILL_41_5_1 gnd vdd FILL
XFILL_78_DFFSR_36 gnd vdd FILL
XFILL_15_DFFSR_169 gnd vdd FILL
XFILL_22_MUX2X1_155 gnd vdd FILL
XFILL_78_DFFSR_47 gnd vdd FILL
XFILL_5_MUX2X1_104 gnd vdd FILL
XFILL_78_DFFSR_58 gnd vdd FILL
XFILL_22_MUX2X1_166 gnd vdd FILL
XFILL_19_DFFSR_102 gnd vdd FILL
XFILL_5_MUX2X1_115 gnd vdd FILL
XFILL_40_0_0 gnd vdd FILL
XFILL_78_DFFSR_69 gnd vdd FILL
XFILL_22_MUX2X1_177 gnd vdd FILL
XFILL_22_MUX2X1_188 gnd vdd FILL
XFILL_19_DFFSR_113 gnd vdd FILL
XFILL_1_INVX1_10 gnd vdd FILL
XFILL_19_DFFSR_124 gnd vdd FILL
XFILL_5_MUX2X1_126 gnd vdd FILL
XFILL_1_INVX1_21 gnd vdd FILL
XFILL_19_DFFSR_135 gnd vdd FILL
XFILL_5_MUX2X1_137 gnd vdd FILL
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XFILL_19_DFFSR_146 gnd vdd FILL
XFILL_1_INVX1_32 gnd vdd FILL
XFILL_5_MUX2X1_148 gnd vdd FILL
XFILL_1_INVX1_43 gnd vdd FILL
XFILL_5_MUX2X1_159 gnd vdd FILL
XFILL_2_AND2X2_2 gnd vdd FILL
XFILL_19_DFFSR_157 gnd vdd FILL
XFILL_1_INVX1_54 gnd vdd FILL
XFILL_1_INVX1_65 gnd vdd FILL
XFILL_19_DFFSR_168 gnd vdd FILL
XFILL_19_DFFSR_179 gnd vdd FILL
XFILL_11_NOR3X1_15 gnd vdd FILL
XFILL_2_OAI22X1_40 gnd vdd FILL
XFILL_47_DFFSR_13 gnd vdd FILL
XFILL_2_OAI22X1_51 gnd vdd FILL
XFILL_1_INVX1_76 gnd vdd FILL
XFILL_11_NOR3X1_26 gnd vdd FILL
XFILL_47_DFFSR_24 gnd vdd FILL
XFILL_1_INVX1_87 gnd vdd FILL
XFILL_47_DFFSR_35 gnd vdd FILL
XFILL_1_INVX1_98 gnd vdd FILL
XFILL_6_OAI21X1_20 gnd vdd FILL
XFILL_11_NOR3X1_37 gnd vdd FILL
XFILL_6_OAI21X1_31 gnd vdd FILL
XFILL_11_NOR3X1_48 gnd vdd FILL
XFILL_61_DFFSR_204 gnd vdd FILL
XFILL_47_DFFSR_46 gnd vdd FILL
XFILL_6_OAI21X1_42 gnd vdd FILL
XFILL_61_DFFSR_215 gnd vdd FILL
XFILL_47_DFFSR_57 gnd vdd FILL
XFILL_47_DFFSR_68 gnd vdd FILL
XFILL_61_DFFSR_226 gnd vdd FILL
XFILL_61_DFFSR_237 gnd vdd FILL
XFILL_47_DFFSR_79 gnd vdd FILL
XFILL_61_DFFSR_248 gnd vdd FILL
XFILL_15_NOR3X1_14 gnd vdd FILL
XFILL_87_DFFSR_12 gnd vdd FILL
XFILL_61_DFFSR_259 gnd vdd FILL
XFILL_87_DFFSR_23 gnd vdd FILL
XFILL_15_NOR3X1_25 gnd vdd FILL
XFILL_15_NOR3X1_36 gnd vdd FILL
XFILL_87_DFFSR_34 gnd vdd FILL
XFILL_15_NOR3X1_47 gnd vdd FILL
XFILL_65_DFFSR_203 gnd vdd FILL
XFILL_87_DFFSR_45 gnd vdd FILL
XFILL_65_DFFSR_214 gnd vdd FILL
XFILL_87_DFFSR_56 gnd vdd FILL
XFILL_16_DFFSR_12 gnd vdd FILL
XFILL_87_DFFSR_67 gnd vdd FILL
XFILL_8_BUFX4_105 gnd vdd FILL
XFILL_16_DFFSR_23 gnd vdd FILL
XFILL_65_DFFSR_225 gnd vdd FILL
XFILL_87_DFFSR_78 gnd vdd FILL
XFILL_65_DFFSR_236 gnd vdd FILL
XFILL_16_DFFSR_34 gnd vdd FILL
XFILL_87_DFFSR_89 gnd vdd FILL
XFILL_65_DFFSR_247 gnd vdd FILL
XFILL_16_DFFSR_45 gnd vdd FILL
XFILL_19_NOR3X1_13 gnd vdd FILL
XFILL_65_DFFSR_258 gnd vdd FILL
XFILL_16_DFFSR_56 gnd vdd FILL
XFILL_19_NOR3X1_24 gnd vdd FILL
XFILL_12_INVX8_4 gnd vdd FILL
XFILL_65_DFFSR_269 gnd vdd FILL
XFILL_16_DFFSR_67 gnd vdd FILL
XFILL_16_DFFSR_78 gnd vdd FILL
XFILL_19_NOR3X1_35 gnd vdd FILL
XFILL_69_DFFSR_202 gnd vdd FILL
XFILL_16_DFFSR_89 gnd vdd FILL
XFILL_19_NOR3X1_46 gnd vdd FILL
XFILL_49_6_1 gnd vdd FILL
XFILL_69_DFFSR_213 gnd vdd FILL
XFILL_60_8 gnd vdd FILL
XFILL_56_DFFSR_11 gnd vdd FILL
XFILL_56_DFFSR_22 gnd vdd FILL
XFILL_69_DFFSR_224 gnd vdd FILL
XFILL_69_DFFSR_235 gnd vdd FILL
XFILL_48_1_0 gnd vdd FILL
XFILL_56_DFFSR_33 gnd vdd FILL
XFILL_27_NOR3X1_8 gnd vdd FILL
XFILL_69_DFFSR_246 gnd vdd FILL
XFILL_56_DFFSR_44 gnd vdd FILL
XFILL_56_DFFSR_55 gnd vdd FILL
XFILL_69_DFFSR_257 gnd vdd FILL
XFILL_69_DFFSR_268 gnd vdd FILL
XFILL_24_CLKBUF1_9 gnd vdd FILL
XFILL_56_DFFSR_66 gnd vdd FILL
XFILL_56_DFFSR_77 gnd vdd FILL
XFILL_56_DFFSR_88 gnd vdd FILL
XFILL_2_NOR2X1_19 gnd vdd FILL
XFILL_56_DFFSR_99 gnd vdd FILL
XFILL_8_NAND3X1_18 gnd vdd FILL
XFILL_8_NAND3X1_29 gnd vdd FILL
XFILL_1_NOR2X1_9 gnd vdd FILL
XFILL_54_DFFSR_4 gnd vdd FILL
XFILL_25_DFFSR_10 gnd vdd FILL
XFILL_25_DFFSR_21 gnd vdd FILL
XFILL_28_CLKBUF1_8 gnd vdd FILL
XFILL_25_DFFSR_32 gnd vdd FILL
XFILL_25_DFFSR_43 gnd vdd FILL
XFILL_6_NOR2X1_18 gnd vdd FILL
XFILL_25_DFFSR_54 gnd vdd FILL
XFILL_32_5_1 gnd vdd FILL
XFILL_6_NOR2X1_29 gnd vdd FILL
XFILL_25_DFFSR_65 gnd vdd FILL
XFILL_25_DFFSR_76 gnd vdd FILL
XFILL_31_0_0 gnd vdd FILL
XFILL_25_DFFSR_87 gnd vdd FILL
XFILL_25_DFFSR_98 gnd vdd FILL
XFILL_65_DFFSR_20 gnd vdd FILL
XFILL_65_DFFSR_31 gnd vdd FILL
XFILL_65_DFFSR_42 gnd vdd FILL
XFILL_0_MUX2X1_7 gnd vdd FILL
XFILL_65_DFFSR_53 gnd vdd FILL
XFILL_65_DFFSR_64 gnd vdd FILL
XFILL_65_DFFSR_75 gnd vdd FILL
XFILL_65_DFFSR_86 gnd vdd FILL
XFILL_15_NAND3X1_105 gnd vdd FILL
XFILL_65_DFFSR_97 gnd vdd FILL
XFILL_6_DFFSR_9 gnd vdd FILL
XFILL_8_DFFSR_11 gnd vdd FILL
XFILL_15_NAND3X1_116 gnd vdd FILL
XFILL_15_NAND3X1_127 gnd vdd FILL
XFILL_8_DFFSR_22 gnd vdd FILL
XFILL_19_DFFSR_7 gnd vdd FILL
XFILL_8_DFFSR_33 gnd vdd FILL
XFILL_8_DFFSR_44 gnd vdd FILL
XFILL_8_DFFSR_55 gnd vdd FILL
XFILL_76_DFFSR_8 gnd vdd FILL
XFILL_34_DFFSR_30 gnd vdd FILL
XFILL_8_DFFSR_66 gnd vdd FILL
XFILL_11_MUX2X1_140 gnd vdd FILL
XFILL_34_DFFSR_41 gnd vdd FILL
XFILL_8_DFFSR_77 gnd vdd FILL
XFILL_34_DFFSR_52 gnd vdd FILL
XFILL_11_MUX2X1_151 gnd vdd FILL
XFILL_34_DFFSR_63 gnd vdd FILL
XFILL_8_DFFSR_88 gnd vdd FILL
XFILL_11_MUX2X1_162 gnd vdd FILL
XFILL_8_DFFSR_99 gnd vdd FILL
XFILL_34_DFFSR_74 gnd vdd FILL
XFILL_11_MUX2X1_173 gnd vdd FILL
XFILL_34_DFFSR_85 gnd vdd FILL
XFILL_81_DFFSR_190 gnd vdd FILL
XFILL_11_MUX2X1_184 gnd vdd FILL
XFILL_34_DFFSR_96 gnd vdd FILL
XFILL_32_DFFSR_203 gnd vdd FILL
XFILL_32_DFFSR_214 gnd vdd FILL
XFILL_74_DFFSR_40 gnd vdd FILL
XFILL_32_DFFSR_225 gnd vdd FILL
XFILL_32_DFFSR_236 gnd vdd FILL
XFILL_74_DFFSR_51 gnd vdd FILL
XFILL_32_DFFSR_247 gnd vdd FILL
XFILL_1_DFFSR_260 gnd vdd FILL
XFILL_32_DFFSR_258 gnd vdd FILL
XFILL_74_DFFSR_62 gnd vdd FILL
XFILL_1_DFFSR_271 gnd vdd FILL
XFILL_74_DFFSR_73 gnd vdd FILL
XFILL_74_DFFSR_84 gnd vdd FILL
XFILL_32_DFFSR_269 gnd vdd FILL
XFILL_74_DFFSR_95 gnd vdd FILL
XFILL_39_1_0 gnd vdd FILL
XFILL_36_DFFSR_202 gnd vdd FILL
XFILL_27_CLKBUF1_19 gnd vdd FILL
XFILL_36_DFFSR_213 gnd vdd FILL
XFILL_36_DFFSR_224 gnd vdd FILL
XFILL_36_DFFSR_235 gnd vdd FILL
XFILL_36_DFFSR_246 gnd vdd FILL
XFILL_5_DFFSR_270 gnd vdd FILL
XFILL_36_DFFSR_257 gnd vdd FILL
XFILL_36_DFFSR_268 gnd vdd FILL
XFILL_14_NOR3X1_3 gnd vdd FILL
XFILL_2_MUX2X1_15 gnd vdd FILL
XFILL_2_MUX2X1_26 gnd vdd FILL
XFILL_43_DFFSR_50 gnd vdd FILL
XFILL_63_DFFSR_102 gnd vdd FILL
XFILL_2_MUX2X1_37 gnd vdd FILL
XFILL_63_DFFSR_113 gnd vdd FILL
XFILL_43_DFFSR_61 gnd vdd FILL
XFILL_63_DFFSR_124 gnd vdd FILL
XFILL_2_MUX2X1_48 gnd vdd FILL
XFILL_43_DFFSR_72 gnd vdd FILL
XFILL_43_DFFSR_83 gnd vdd FILL
XFILL_63_DFFSR_135 gnd vdd FILL
XFILL_2_MUX2X1_59 gnd vdd FILL
XFILL_63_DFFSR_146 gnd vdd FILL
XFILL_10_NAND3X1_101 gnd vdd FILL
XFILL_43_DFFSR_94 gnd vdd FILL
XFILL_63_DFFSR_157 gnd vdd FILL
XFILL_10_NAND3X1_112 gnd vdd FILL
XFILL_63_DFFSR_168 gnd vdd FILL
XFILL_10_NAND3X1_123 gnd vdd FILL
XFILL_23_5_1 gnd vdd FILL
XFILL_63_DFFSR_179 gnd vdd FILL
XFILL_6_MUX2X1_14 gnd vdd FILL
XFILL_6_MUX2X1_25 gnd vdd FILL
XFILL_67_DFFSR_101 gnd vdd FILL
XFILL_22_0_0 gnd vdd FILL
XFILL_83_DFFSR_60 gnd vdd FILL
XFILL_6_MUX2X1_36 gnd vdd FILL
XFILL_6_MUX2X1_47 gnd vdd FILL
XFILL_67_DFFSR_112 gnd vdd FILL
XFILL_8_NOR2X1_108 gnd vdd FILL
XFILL_83_DFFSR_71 gnd vdd FILL
XFILL_67_DFFSR_123 gnd vdd FILL
XFILL_83_DFFSR_82 gnd vdd FILL
XFILL_67_DFFSR_134 gnd vdd FILL
XFILL_6_MUX2X1_58 gnd vdd FILL
XFILL_8_NOR2X1_119 gnd vdd FILL
XFILL_6_MUX2X1_69 gnd vdd FILL
XFILL_83_DFFSR_93 gnd vdd FILL
XFILL_67_DFFSR_145 gnd vdd FILL
XFILL_14_NAND3X1_10 gnd vdd FILL
XFILL_10_OAI21X1_2 gnd vdd FILL
XFILL_14_NAND3X1_21 gnd vdd FILL
XFILL_12_DFFSR_60 gnd vdd FILL
XFILL_67_DFFSR_156 gnd vdd FILL
XFILL_0_BUFX4_9 gnd vdd FILL
XFILL_67_DFFSR_167 gnd vdd FILL
XFILL_14_NAND3X1_32 gnd vdd FILL
XFILL_12_DFFSR_71 gnd vdd FILL
XFILL_12_DFFSR_82 gnd vdd FILL
XFILL_67_DFFSR_178 gnd vdd FILL
XFILL_1_MUX2X1_190 gnd vdd FILL
XFILL_14_NAND3X1_43 gnd vdd FILL
XFILL_13_BUFX4_7 gnd vdd FILL
XFILL_12_DFFSR_93 gnd vdd FILL
XFILL_67_DFFSR_189 gnd vdd FILL
XFILL_14_NAND3X1_54 gnd vdd FILL
XFILL_14_NAND3X1_65 gnd vdd FILL
XFILL_34_CLKBUF1_10 gnd vdd FILL
XFILL_34_CLKBUF1_21 gnd vdd FILL
XFILL_14_NAND3X1_76 gnd vdd FILL
XFILL_23_NOR3X1_1 gnd vdd FILL
XFILL_34_CLKBUF1_32 gnd vdd FILL
XFILL_14_NAND3X1_87 gnd vdd FILL
XFILL_14_OAI21X1_1 gnd vdd FILL
XFILL_14_NAND3X1_98 gnd vdd FILL
XFILL_1_NAND3X1_106 gnd vdd FILL
XFILL_1_NAND3X1_117 gnd vdd FILL
XFILL_52_DFFSR_70 gnd vdd FILL
XFILL_1_NAND3X1_128 gnd vdd FILL
XFILL_52_DFFSR_81 gnd vdd FILL
XFILL_52_DFFSR_92 gnd vdd FILL
XFILL_11_NOR2X1_70 gnd vdd FILL
XFILL_11_NOR2X1_81 gnd vdd FILL
XFILL_11_NOR2X1_92 gnd vdd FILL
XFILL_22_MUX2X1_12 gnd vdd FILL
XFILL_22_MUX2X1_23 gnd vdd FILL
XFILL_21_DFFSR_80 gnd vdd FILL
XFILL_22_MUX2X1_34 gnd vdd FILL
XFILL_22_MUX2X1_45 gnd vdd FILL
XFILL_6_6_1 gnd vdd FILL
XFILL_21_DFFSR_91 gnd vdd FILL
XFILL_6_NOR3X1_2 gnd vdd FILL
XFILL_22_MUX2X1_56 gnd vdd FILL
XFILL_5_OAI22X1_17 gnd vdd FILL
XFILL_5_1_0 gnd vdd FILL
XFILL_22_MUX2X1_67 gnd vdd FILL
XFILL_22_MUX2X1_78 gnd vdd FILL
XFILL_5_OAI22X1_28 gnd vdd FILL
XFILL_22_MUX2X1_89 gnd vdd FILL
XFILL_5_OAI22X1_39 gnd vdd FILL
XFILL_18_AOI22X1_10 gnd vdd FILL
XFILL_9_OAI21X1_19 gnd vdd FILL
XFILL_61_DFFSR_90 gnd vdd FILL
XFILL_4_NAND3X1_60 gnd vdd FILL
XFILL_4_NAND3X1_71 gnd vdd FILL
XFILL_4_NAND3X1_82 gnd vdd FILL
XFILL_36_DFFSR_1 gnd vdd FILL
XFILL_4_NAND3X1_93 gnd vdd FILL
XFILL_30_DFFSR_102 gnd vdd FILL
XFILL_8_NAND2X1_40 gnd vdd FILL
XFILL_8_NAND2X1_51 gnd vdd FILL
XFILL_30_DFFSR_113 gnd vdd FILL
XFILL_30_DFFSR_124 gnd vdd FILL
XFILL_8_NAND2X1_62 gnd vdd FILL
XFILL_4_DFFSR_70 gnd vdd FILL
XFILL_14_5_1 gnd vdd FILL
XFILL_8_NAND2X1_73 gnd vdd FILL
XFILL_30_DFFSR_135 gnd vdd FILL
XFILL_4_DFFSR_81 gnd vdd FILL
XFILL_30_DFFSR_146 gnd vdd FILL
XFILL_4_DFFSR_92 gnd vdd FILL
XFILL_13_0_0 gnd vdd FILL
XFILL_8_NAND2X1_84 gnd vdd FILL
XFILL_30_DFFSR_157 gnd vdd FILL
XFILL_8_NAND2X1_95 gnd vdd FILL
XFILL_30_DFFSR_168 gnd vdd FILL
XFILL_30_DFFSR_179 gnd vdd FILL
XFILL_34_DFFSR_101 gnd vdd FILL
XFILL_11_NAND2X1_3 gnd vdd FILL
XFILL_16_CLKBUF1_15 gnd vdd FILL
XFILL_34_DFFSR_112 gnd vdd FILL
XFILL_16_CLKBUF1_26 gnd vdd FILL
XFILL_34_DFFSR_123 gnd vdd FILL
XFILL_34_DFFSR_134 gnd vdd FILL
XFILL_16_CLKBUF1_37 gnd vdd FILL
XFILL_34_DFFSR_145 gnd vdd FILL
XFILL_11_AOI21X1_12 gnd vdd FILL
XFILL_34_DFFSR_156 gnd vdd FILL
XFILL_11_AOI21X1_23 gnd vdd FILL
XFILL_11_AOI21X1_34 gnd vdd FILL
XFILL_3_DFFSR_180 gnd vdd FILL
XFILL_34_DFFSR_167 gnd vdd FILL
XFILL_11_AOI21X1_45 gnd vdd FILL
XFILL_34_DFFSR_178 gnd vdd FILL
XFILL_3_DFFSR_191 gnd vdd FILL
XFILL_38_DFFSR_100 gnd vdd FILL
XFILL_34_DFFSR_189 gnd vdd FILL
XAND2X2_3 AND2X2_6/A AND2X2_3/B gnd AND2X2_3/Y vdd AND2X2
XFILL_11_AOI21X1_56 gnd vdd FILL
XFILL_20_DFFSR_7 gnd vdd FILL
XFILL_11_AOI21X1_67 gnd vdd FILL
XFILL_38_DFFSR_111 gnd vdd FILL
XFILL_11_AOI21X1_78 gnd vdd FILL
XFILL_38_DFFSR_122 gnd vdd FILL
XFILL_38_DFFSR_133 gnd vdd FILL
XFILL_38_DFFSR_144 gnd vdd FILL
XFILL_38_DFFSR_155 gnd vdd FILL
XFILL_58_DFFSR_5 gnd vdd FILL
XFILL_38_DFFSR_166 gnd vdd FILL
XFILL_38_DFFSR_177 gnd vdd FILL
XFILL_30_NOR3X1_13 gnd vdd FILL
XFILL_7_DFFSR_190 gnd vdd FILL
XFILL_38_DFFSR_188 gnd vdd FILL
XFILL_30_NOR3X1_24 gnd vdd FILL
XFILL_38_DFFSR_199 gnd vdd FILL
XFILL_30_NOR3X1_35 gnd vdd FILL
XFILL_80_DFFSR_202 gnd vdd FILL
XFILL_30_NOR3X1_46 gnd vdd FILL
XFILL_80_DFFSR_213 gnd vdd FILL
XFILL_2_3 gnd vdd FILL
XFILL_80_DFFSR_224 gnd vdd FILL
XFILL_80_DFFSR_235 gnd vdd FILL
XFILL_80_DFFSR_246 gnd vdd FILL
XFILL_80_DFFSR_257 gnd vdd FILL
XFILL_80_DFFSR_268 gnd vdd FILL
XFILL_84_DFFSR_201 gnd vdd FILL
XFILL_84_DFFSR_212 gnd vdd FILL
XFILL_84_DFFSR_223 gnd vdd FILL
XFILL_84_DFFSR_234 gnd vdd FILL
XFILL_11_AOI21X1_8 gnd vdd FILL
XFILL_0_BUFX4_19 gnd vdd FILL
XFILL_84_DFFSR_245 gnd vdd FILL
XFILL_64_4_1 gnd vdd FILL
XFILL_6_CLKBUF1_10 gnd vdd FILL
XFILL_84_DFFSR_256 gnd vdd FILL
XFILL_6_CLKBUF1_21 gnd vdd FILL
XFILL_84_DFFSR_267 gnd vdd FILL
XFILL_44_3 gnd vdd FILL
XFILL_6_CLKBUF1_32 gnd vdd FILL
XFILL_14_MUX2X1_106 gnd vdd FILL
XFILL_0_INVX1_140 gnd vdd FILL
XFILL_14_MUX2X1_117 gnd vdd FILL
XFILL_15_AOI21X1_7 gnd vdd FILL
XFILL_0_INVX1_151 gnd vdd FILL
XFILL_14_MUX2X1_128 gnd vdd FILL
XFILL_0_INVX1_162 gnd vdd FILL
XFILL_1_AOI21X1_40 gnd vdd FILL
XFILL_14_MUX2X1_139 gnd vdd FILL
XFILL_1_AOI21X1_51 gnd vdd FILL
XFILL_0_INVX1_173 gnd vdd FILL
XFILL_0_INVX1_184 gnd vdd FILL
XFILL_1_AOI21X1_62 gnd vdd FILL
XFILL_11_OAI22X1_20 gnd vdd FILL
XFILL_0_INVX1_195 gnd vdd FILL
XFILL_11_OAI22X1_31 gnd vdd FILL
XFILL_1_AOI21X1_73 gnd vdd FILL
XFILL_11_OAI22X1_42 gnd vdd FILL
XFILL_15_OAI21X1_11 gnd vdd FILL
XFILL_4_INVX1_150 gnd vdd FILL
XFILL_15_OAI21X1_22 gnd vdd FILL
XFILL_4_INVX1_161 gnd vdd FILL
XFILL_15_OAI21X1_33 gnd vdd FILL
XFILL_4_NOR2X1_150 gnd vdd FILL
XFILL_15_OAI21X1_44 gnd vdd FILL
XFILL_4_INVX1_172 gnd vdd FILL
XFILL_4_INVX1_183 gnd vdd FILL
XFILL_4_NOR2X1_161 gnd vdd FILL
XFILL_4_INVX1_194 gnd vdd FILL
XFILL_4_NOR2X1_172 gnd vdd FILL
XFILL_4_NOR2X1_183 gnd vdd FILL
XFILL_4_NOR2X1_194 gnd vdd FILL
XFILL_2_OAI22X1_1 gnd vdd FILL
XFILL_21_MUX2X1_130 gnd vdd FILL
XFILL_21_MUX2X1_141 gnd vdd FILL
XFILL_21_MUX2X1_152 gnd vdd FILL
XFILL_21_MUX2X1_163 gnd vdd FILL
XFILL_60_11 gnd vdd FILL
XFILL_4_MUX2X1_101 gnd vdd FILL
XFILL_4_MUX2X1_112 gnd vdd FILL
XFILL_21_MUX2X1_174 gnd vdd FILL
XNAND3X1_19 INVX1_164/A BUFX4_90/Y NOR3X1_51/Y gnd OAI21X1_27/C vdd NAND3X1
XFILL_21_MUX2X1_185 gnd vdd FILL
XFILL_4_MUX2X1_123 gnd vdd FILL
XFILL_4_MUX2X1_134 gnd vdd FILL
XFILL_4_MUX2X1_145 gnd vdd FILL
XFILL_4_MUX2X1_156 gnd vdd FILL
XFILL_4_MUX2X1_167 gnd vdd FILL
XFILL_35_DFFSR_19 gnd vdd FILL
XFILL_4_MUX2X1_178 gnd vdd FILL
XFILL_4_MUX2X1_189 gnd vdd FILL
XNOR2X1_19 NOR2X1_19/A NOR2X1_19/B gnd NOR2X1_19/Y vdd NOR2X1
XFILL_51_DFFSR_201 gnd vdd FILL
XFILL_55_4_1 gnd vdd FILL
XFILL_51_DFFSR_212 gnd vdd FILL
XFILL_5_OAI21X1_50 gnd vdd FILL
XFILL_51_DFFSR_223 gnd vdd FILL
XFILL_51_DFFSR_234 gnd vdd FILL
XFILL_51_DFFSR_245 gnd vdd FILL
XFILL_75_DFFSR_18 gnd vdd FILL
XFILL_51_DFFSR_256 gnd vdd FILL
XFILL_75_DFFSR_29 gnd vdd FILL
XFILL_51_DFFSR_267 gnd vdd FILL
XFILL_55_DFFSR_200 gnd vdd FILL
XFILL_18_MUX2X1_8 gnd vdd FILL
XFILL_55_DFFSR_211 gnd vdd FILL
XFILL_55_DFFSR_222 gnd vdd FILL
XFILL_55_DFFSR_233 gnd vdd FILL
XFILL_11_NAND3X1_102 gnd vdd FILL
XFILL_11_NAND3X1_113 gnd vdd FILL
XFILL_55_DFFSR_244 gnd vdd FILL
XFILL_55_DFFSR_255 gnd vdd FILL
XFILL_9_BUFX4_30 gnd vdd FILL
XFILL_11_NAND3X1_124 gnd vdd FILL
XFILL_55_DFFSR_266 gnd vdd FILL
XFILL_10_CLKBUF1_7 gnd vdd FILL
XFILL_9_BUFX4_41 gnd vdd FILL
XFILL_9_BUFX4_52 gnd vdd FILL
XFILL_82_DFFSR_100 gnd vdd FILL
XFILL_9_BUFX4_63 gnd vdd FILL
XFILL_59_DFFSR_210 gnd vdd FILL
XFILL_44_DFFSR_17 gnd vdd FILL
XFILL_82_DFFSR_111 gnd vdd FILL
XFILL_0_BUFX2_6 gnd vdd FILL
XFILL_44_DFFSR_28 gnd vdd FILL
XFILL_59_DFFSR_221 gnd vdd FILL
XFILL_9_BUFX4_74 gnd vdd FILL
XFILL_82_DFFSR_122 gnd vdd FILL
XFILL_82_DFFSR_133 gnd vdd FILL
XFILL_9_BUFX4_85 gnd vdd FILL
XFILL_44_DFFSR_39 gnd vdd FILL
XFILL_9_BUFX4_96 gnd vdd FILL
XFILL_82_DFFSR_144 gnd vdd FILL
XFILL_59_DFFSR_232 gnd vdd FILL
XFILL_59_DFFSR_243 gnd vdd FILL
XFILL_82_DFFSR_155 gnd vdd FILL
XFILL_59_DFFSR_254 gnd vdd FILL
XFILL_82_DFFSR_166 gnd vdd FILL
XFILL_59_DFFSR_265 gnd vdd FILL
XFILL_82_DFFSR_177 gnd vdd FILL
XFILL_14_CLKBUF1_6 gnd vdd FILL
XFILL_82_DFFSR_188 gnd vdd FILL
XFILL_2_DFFSR_203 gnd vdd FILL
XFILL_82_DFFSR_199 gnd vdd FILL
XFILL_2_DFFSR_214 gnd vdd FILL
XFILL_84_DFFSR_16 gnd vdd FILL
XFILL_86_DFFSR_110 gnd vdd FILL
XFILL_7_NAND3X1_15 gnd vdd FILL
XFILL_84_DFFSR_27 gnd vdd FILL
XFILL_86_DFFSR_121 gnd vdd FILL
XFILL_2_DFFSR_225 gnd vdd FILL
XFILL_86_DFFSR_132 gnd vdd FILL
XFILL_7_NAND3X1_26 gnd vdd FILL
XFILL_84_DFFSR_38 gnd vdd FILL
XFILL_2_DFFSR_236 gnd vdd FILL
XFILL_86_DFFSR_143 gnd vdd FILL
XFILL_2_DFFSR_247 gnd vdd FILL
XFILL_84_DFFSR_49 gnd vdd FILL
XFILL_7_NAND3X1_37 gnd vdd FILL
XFILL_86_DFFSR_154 gnd vdd FILL
XFILL_2_NAND3X1_107 gnd vdd FILL
XFILL_2_DFFSR_258 gnd vdd FILL
XFILL_10_BUFX4_101 gnd vdd FILL
XFILL_2_NAND3X1_118 gnd vdd FILL
XFILL_13_DFFSR_16 gnd vdd FILL
XFILL_7_NAND3X1_48 gnd vdd FILL
XFILL_7_NAND3X1_59 gnd vdd FILL
XFILL_2_DFFSR_269 gnd vdd FILL
XFILL_2_NAND3X1_129 gnd vdd FILL
XFILL_86_DFFSR_165 gnd vdd FILL
XFILL_13_DFFSR_27 gnd vdd FILL
XFILL_13_DFFSR_38 gnd vdd FILL
XFILL_86_DFFSR_176 gnd vdd FILL
XFILL_18_CLKBUF1_5 gnd vdd FILL
XFILL_6_DFFSR_202 gnd vdd FILL
XFILL_86_DFFSR_187 gnd vdd FILL
XFILL_13_DFFSR_49 gnd vdd FILL
XFILL_6_DFFSR_213 gnd vdd FILL
XFILL_86_DFFSR_198 gnd vdd FILL
XFILL_3_NAND3X1_2 gnd vdd FILL
XFILL_6_DFFSR_224 gnd vdd FILL
XFILL_6_DFFSR_235 gnd vdd FILL
XFILL_6_DFFSR_246 gnd vdd FILL
XFILL_6_DFFSR_257 gnd vdd FILL
XFILL_14_BUFX4_100 gnd vdd FILL
XFILL_6_DFFSR_268 gnd vdd FILL
XFILL_53_DFFSR_15 gnd vdd FILL
XFILL_53_DFFSR_26 gnd vdd FILL
XFILL_53_DFFSR_37 gnd vdd FILL
XFILL_53_DFFSR_48 gnd vdd FILL
XFILL_7_NAND3X1_1 gnd vdd FILL
XFILL_53_DFFSR_59 gnd vdd FILL
XMUX2X1_15 BUFX4_83/Y INVX1_28/Y MUX2X1_16/S gnd DFFSR_23/D vdd MUX2X1
XFILL_0_NAND2X1_17 gnd vdd FILL
XFILL_46_4_1 gnd vdd FILL
XFILL_0_NAND2X1_28 gnd vdd FILL
XMUX2X1_26 BUFX4_63/Y INVX1_39/Y NOR2X1_12/B gnd MUX2X1_26/Y vdd MUX2X1
XMUX2X1_37 INVX1_50/Y BUFX4_86/Y NAND2X1_5/Y gnd MUX2X1_37/Y vdd MUX2X1
XFILL_0_NAND2X1_39 gnd vdd FILL
XFILL_24_DFFSR_8 gnd vdd FILL
XMUX2X1_48 INVX1_61/Y BUFX4_77/Y NAND2X1_7/Y gnd MUX2X1_48/Y vdd MUX2X1
XFILL_22_DFFSR_14 gnd vdd FILL
XNOR2X1_109 INVX2_4/A INVX2_5/A gnd INVX1_57/A vdd NOR2X1
XMUX2X1_59 BUFX4_85/Y INVX1_72/Y NOR2X1_22/Y gnd MUX2X1_59/Y vdd MUX2X1
XFILL_81_DFFSR_9 gnd vdd FILL
XFILL_22_DFFSR_25 gnd vdd FILL
XFILL_22_DFFSR_36 gnd vdd FILL
XFILL_22_DFFSR_47 gnd vdd FILL
XFILL_22_DFFSR_58 gnd vdd FILL
XFILL_13_BUFX4_90 gnd vdd FILL
XFILL_22_DFFSR_69 gnd vdd FILL
XFILL_10_MUX2X1_170 gnd vdd FILL
XFILL_62_DFFSR_13 gnd vdd FILL
XFILL_23_8 gnd vdd FILL
XFILL_10_MUX2X1_181 gnd vdd FILL
XFILL_22_DFFSR_200 gnd vdd FILL
XFILL_62_DFFSR_24 gnd vdd FILL
XFILL_10_MUX2X1_192 gnd vdd FILL
XFILL_22_DFFSR_211 gnd vdd FILL
XFILL_62_DFFSR_35 gnd vdd FILL
XFILL_22_DFFSR_222 gnd vdd FILL
XFILL_62_DFFSR_46 gnd vdd FILL
XFILL_16_7 gnd vdd FILL
XFILL_3_AOI22X1_7 gnd vdd FILL
XFILL_62_DFFSR_57 gnd vdd FILL
XFILL_22_DFFSR_233 gnd vdd FILL
XFILL_62_DFFSR_68 gnd vdd FILL
XFILL_22_DFFSR_244 gnd vdd FILL
XFILL_22_DFFSR_255 gnd vdd FILL
XFILL_62_DFFSR_79 gnd vdd FILL
XFILL_22_DFFSR_266 gnd vdd FILL
XFILL_3_INVX1_206 gnd vdd FILL
XFILL_26_DFFSR_210 gnd vdd FILL
XFILL_26_CLKBUF1_16 gnd vdd FILL
XFILL_3_INVX1_217 gnd vdd FILL
XFILL_5_DFFSR_15 gnd vdd FILL
XFILL_26_DFFSR_221 gnd vdd FILL
XFILL_3_INVX1_228 gnd vdd FILL
XDFFSR_7 DFFSR_7/Q DFFSR_7/CLK DFFSR_8/R vdd DFFSR_7/D gnd vdd DFFSR
XFILL_26_CLKBUF1_27 gnd vdd FILL
XFILL_26_CLKBUF1_38 gnd vdd FILL
XFILL_7_AOI22X1_6 gnd vdd FILL
XFILL_5_DFFSR_26 gnd vdd FILL
XFILL_31_DFFSR_12 gnd vdd FILL
XFILL_5_DFFSR_37 gnd vdd FILL
XFILL_26_DFFSR_232 gnd vdd FILL
XFILL_26_DFFSR_243 gnd vdd FILL
XFILL_5_DFFSR_48 gnd vdd FILL
XFILL_31_DFFSR_23 gnd vdd FILL
XFILL_26_DFFSR_254 gnd vdd FILL
XFILL_31_DFFSR_34 gnd vdd FILL
XFILL_5_DFFSR_59 gnd vdd FILL
XFILL_26_DFFSR_265 gnd vdd FILL
XFILL_31_DFFSR_45 gnd vdd FILL
XFILL_31_DFFSR_56 gnd vdd FILL
XFILL_7_INVX1_205 gnd vdd FILL
XFILL_31_DFFSR_67 gnd vdd FILL
XFILL_7_INVX1_216 gnd vdd FILL
XFILL_31_DFFSR_78 gnd vdd FILL
XFILL_53_DFFSR_110 gnd vdd FILL
XFILL_31_DFFSR_89 gnd vdd FILL
XFILL_7_INVX1_80 gnd vdd FILL
XFILL_4_AOI21X1_17 gnd vdd FILL
XFILL_7_INVX1_227 gnd vdd FILL
XFILL_53_DFFSR_121 gnd vdd FILL
XFILL_53_DFFSR_132 gnd vdd FILL
XFILL_7_INVX1_91 gnd vdd FILL
XFILL_53_DFFSR_143 gnd vdd FILL
XFILL_71_DFFSR_11 gnd vdd FILL
XFILL_4_AOI21X1_28 gnd vdd FILL
XFILL_4_AOI21X1_39 gnd vdd FILL
XFILL_71_DFFSR_22 gnd vdd FILL
XFILL_53_DFFSR_154 gnd vdd FILL
XFILL_71_DFFSR_33 gnd vdd FILL
XFILL_53_DFFSR_165 gnd vdd FILL
XFILL_71_DFFSR_44 gnd vdd FILL
XFILL_14_MUX2X1_1 gnd vdd FILL
XFILL_14_OAI22X1_19 gnd vdd FILL
XFILL_53_DFFSR_176 gnd vdd FILL
XFILL_71_DFFSR_55 gnd vdd FILL
XFILL_53_DFFSR_187 gnd vdd FILL
XFILL_53_DFFSR_198 gnd vdd FILL
XFILL_71_DFFSR_66 gnd vdd FILL
XFILL_71_DFFSR_77 gnd vdd FILL
XFILL_7_NOR2X1_105 gnd vdd FILL
XFILL_57_DFFSR_120 gnd vdd FILL
XFILL_71_DFFSR_88 gnd vdd FILL
XFILL_57_DFFSR_131 gnd vdd FILL
XFILL_71_DFFSR_99 gnd vdd FILL
XFILL_7_NOR2X1_116 gnd vdd FILL
XFILL_57_DFFSR_142 gnd vdd FILL
XFILL_7_NOR2X1_127 gnd vdd FILL
XFILL_57_DFFSR_153 gnd vdd FILL
XFILL_7_NOR2X1_138 gnd vdd FILL
XFILL_7_NOR2X1_149 gnd vdd FILL
XFILL_57_DFFSR_164 gnd vdd FILL
XNAND2X1_30 BUFX4_104/Y NOR3X1_51/Y gnd OAI22X1_9/B vdd NAND2X1
XFILL_57_DFFSR_175 gnd vdd FILL
XNAND2X1_41 NOR2X1_11/A NOR2X1_50/Y gnd NAND3X1_53/A vdd NAND2X1
XFILL_13_NAND3X1_40 gnd vdd FILL
XFILL_0_DFFSR_102 gnd vdd FILL
XNAND2X1_52 BUFX4_88/Y NOR2X1_29/Y gnd OAI22X1_4/D vdd NAND2X1
XFILL_57_DFFSR_186 gnd vdd FILL
XFILL_40_DFFSR_10 gnd vdd FILL
XFILL_13_NAND3X1_51 gnd vdd FILL
XFILL_13_NAND3X1_62 gnd vdd FILL
XFILL_40_DFFSR_21 gnd vdd FILL
XFILL_57_DFFSR_197 gnd vdd FILL
XNAND2X1_63 INVX1_64/A NOR2X1_69/Y gnd NAND3X1_90/A vdd NAND2X1
XFILL_0_DFFSR_113 gnd vdd FILL
XFILL_0_DFFSR_124 gnd vdd FILL
XFILL_13_NAND3X1_73 gnd vdd FILL
XFILL_40_DFFSR_32 gnd vdd FILL
XFILL_40_DFFSR_43 gnd vdd FILL
XNAND2X1_74 NOR2X1_95/Y NOR2X1_94/Y gnd NOR3X1_35/B vdd NAND2X1
XFILL_0_DFFSR_135 gnd vdd FILL
XFILL_11_NOR3X1_7 gnd vdd FILL
XFILL_0_DFFSR_146 gnd vdd FILL
XFILL_13_NAND3X1_84 gnd vdd FILL
XFILL_37_4_1 gnd vdd FILL
XNAND2X1_85 AND2X2_7/A INVX1_57/A gnd NOR2X1_20/A vdd NAND2X1
XFILL_40_DFFSR_54 gnd vdd FILL
XFILL_13_NAND3X1_95 gnd vdd FILL
XFILL_33_CLKBUF1_40 gnd vdd FILL
XNAND2X1_96 OAI21X1_46/B NOR2X1_138/A gnd NAND3X1_37/C vdd NAND2X1
XFILL_0_DFFSR_157 gnd vdd FILL
XFILL_40_DFFSR_65 gnd vdd FILL
XFILL_40_DFFSR_76 gnd vdd FILL
XFILL_0_DFFSR_168 gnd vdd FILL
XFILL_0_DFFSR_179 gnd vdd FILL
XFILL_40_DFFSR_87 gnd vdd FILL
XFILL_40_DFFSR_98 gnd vdd FILL
XFILL_4_DFFSR_101 gnd vdd FILL
XFILL_80_DFFSR_20 gnd vdd FILL
XFILL_4_DFFSR_112 gnd vdd FILL
XFILL_80_DFFSR_31 gnd vdd FILL
XFILL_4_DFFSR_123 gnd vdd FILL
XFILL_4_DFFSR_134 gnd vdd FILL
XFILL_80_DFFSR_42 gnd vdd FILL
XFILL_4_DFFSR_145 gnd vdd FILL
XFILL_80_DFFSR_53 gnd vdd FILL
XFILL_80_DFFSR_64 gnd vdd FILL
XFILL_4_DFFSR_156 gnd vdd FILL
XFILL_4_DFFSR_167 gnd vdd FILL
XFILL_80_DFFSR_75 gnd vdd FILL
XFILL_4_DFFSR_178 gnd vdd FILL
XFILL_80_DFFSR_86 gnd vdd FILL
XFILL_8_DFFSR_100 gnd vdd FILL
XFILL_4_DFFSR_189 gnd vdd FILL
XFILL_80_DFFSR_97 gnd vdd FILL
XFILL_8_DFFSR_111 gnd vdd FILL
XFILL_7_NOR2X1_2 gnd vdd FILL
XFILL_39_DFFSR_109 gnd vdd FILL
XFILL_8_DFFSR_122 gnd vdd FILL
XFILL_12_MUX2X1_20 gnd vdd FILL
XFILL_8_DFFSR_133 gnd vdd FILL
XFILL_12_MUX2X1_31 gnd vdd FILL
XFILL_8_DFFSR_144 gnd vdd FILL
XFILL_12_MUX2X1_42 gnd vdd FILL
XFILL_20_3_1 gnd vdd FILL
XFILL_12_MUX2X1_53 gnd vdd FILL
XFILL_8_DFFSR_155 gnd vdd FILL
XFILL_4_OAI22X1_14 gnd vdd FILL
XFILL_12_MUX2X1_64 gnd vdd FILL
XFILL_8_DFFSR_166 gnd vdd FILL
XFILL_8_DFFSR_177 gnd vdd FILL
XFILL_0_NOR3X1_13 gnd vdd FILL
XFILL_12_MUX2X1_75 gnd vdd FILL
XFILL_4_OAI22X1_25 gnd vdd FILL
XFILL_20_NOR3X1_5 gnd vdd FILL
XFILL_12_MUX2X1_86 gnd vdd FILL
XFILL_0_NOR3X1_24 gnd vdd FILL
XFILL_8_DFFSR_188 gnd vdd FILL
XFILL_4_OAI22X1_36 gnd vdd FILL
XFILL_12_MUX2X1_97 gnd vdd FILL
XFILL_4_OAI22X1_47 gnd vdd FILL
XFILL_8_DFFSR_199 gnd vdd FILL
XFILL_0_NOR3X1_35 gnd vdd FILL
XFILL_0_NOR3X1_46 gnd vdd FILL
XFILL_8_OAI21X1_16 gnd vdd FILL
XFILL_8_OAI21X1_27 gnd vdd FILL
XFILL_16_MUX2X1_30 gnd vdd FILL
XFILL_8_OAI21X1_38 gnd vdd FILL
XFILL_16_MUX2X1_41 gnd vdd FILL
XFILL_16_MUX2X1_52 gnd vdd FILL
XFILL_8_OAI21X1_49 gnd vdd FILL
XFILL_16_MUX2X1_63 gnd vdd FILL
XFILL_4_NOR3X1_12 gnd vdd FILL
XFILL_16_MUX2X1_74 gnd vdd FILL
XFILL_16_MUX2X1_85 gnd vdd FILL
XFILL_4_NOR3X1_23 gnd vdd FILL
XFILL_16_MUX2X1_96 gnd vdd FILL
XFILL_41_DFFSR_2 gnd vdd FILL
XFILL_4_NOR3X1_34 gnd vdd FILL
XFILL_9_DFFSR_1 gnd vdd FILL
XFILL_4_NOR3X1_45 gnd vdd FILL
XFILL_3_NAND3X1_90 gnd vdd FILL
XFILL_20_DFFSR_110 gnd vdd FILL
XFILL_1_NOR2X1_205 gnd vdd FILL
XFILL_20_DFFSR_121 gnd vdd FILL
XFILL_20_DFFSR_132 gnd vdd FILL
XFILL_7_NAND2X1_70 gnd vdd FILL
XFILL_20_DFFSR_143 gnd vdd FILL
XFILL_7_NAND2X1_81 gnd vdd FILL
XFILL_20_DFFSR_154 gnd vdd FILL
XFILL_8_NOR3X1_11 gnd vdd FILL
XFILL_7_NAND2X1_92 gnd vdd FILL
XFILL_20_DFFSR_165 gnd vdd FILL
XFILL_8_NOR3X1_22 gnd vdd FILL
XFILL_8_NOR3X1_33 gnd vdd FILL
XFILL_3_NOR3X1_6 gnd vdd FILL
XFILL_20_DFFSR_176 gnd vdd FILL
XFILL_1_INVX1_105 gnd vdd FILL
XFILL_20_DFFSR_187 gnd vdd FILL
XFILL_20_DFFSR_198 gnd vdd FILL
XFILL_1_INVX1_116 gnd vdd FILL
XFILL_8_NOR3X1_44 gnd vdd FILL
XFILL_15_CLKBUF1_12 gnd vdd FILL
XFILL_1_INVX1_127 gnd vdd FILL
XFILL_4_BUFX2_7 gnd vdd FILL
XFILL_24_DFFSR_120 gnd vdd FILL
XFILL_15_CLKBUF1_23 gnd vdd FILL
XFILL_1_INVX1_138 gnd vdd FILL
XFILL_24_DFFSR_131 gnd vdd FILL
XFILL_15_CLKBUF1_34 gnd vdd FILL
XFILL_24_DFFSR_142 gnd vdd FILL
XFILL_1_INVX1_149 gnd vdd FILL
XFILL_24_DFFSR_153 gnd vdd FILL
XFILL_10_AOI21X1_20 gnd vdd FILL
XFILL_10_AOI21X1_31 gnd vdd FILL
XFILL_24_DFFSR_164 gnd vdd FILL
XFILL_5_INVX1_104 gnd vdd FILL
XFILL_10_AOI21X1_42 gnd vdd FILL
XFILL_24_DFFSR_175 gnd vdd FILL
XFILL_28_4_1 gnd vdd FILL
XFILL_24_DFFSR_186 gnd vdd FILL
XFILL_3_4_1 gnd vdd FILL
XFILL_10_AOI21X1_53 gnd vdd FILL
XFILL_5_INVX1_115 gnd vdd FILL
XFILL_24_DFFSR_197 gnd vdd FILL
XFILL_5_INVX1_126 gnd vdd FILL
XFILL_1_DFFSR_30 gnd vdd FILL
XFILL_10_AOI21X1_64 gnd vdd FILL
XFILL_5_INVX1_137 gnd vdd FILL
XFILL_10_AOI21X1_75 gnd vdd FILL
XFILL_28_DFFSR_130 gnd vdd FILL
XFILL_1_DFFSR_41 gnd vdd FILL
XFILL_5_INVX1_148 gnd vdd FILL
XFILL_1_DFFSR_52 gnd vdd FILL
XFILL_28_DFFSR_141 gnd vdd FILL
XFILL_5_INVX1_159 gnd vdd FILL
XFILL_1_DFFSR_63 gnd vdd FILL
XFILL_28_DFFSR_152 gnd vdd FILL
XFILL_63_DFFSR_6 gnd vdd FILL
XFILL_1_DFFSR_74 gnd vdd FILL
XFILL_28_DFFSR_163 gnd vdd FILL
XFILL_1_DFFSR_85 gnd vdd FILL
XFILL_28_DFFSR_174 gnd vdd FILL
XFILL_20_NOR3X1_10 gnd vdd FILL
XFILL_1_DFFSR_96 gnd vdd FILL
XFILL_28_DFFSR_185 gnd vdd FILL
XFILL_20_NOR3X1_21 gnd vdd FILL
XFILL_28_DFFSR_196 gnd vdd FILL
XFILL_20_NOR3X1_32 gnd vdd FILL
XFILL_15_OR2X2_1 gnd vdd FILL
XFILL_20_NOR3X1_43 gnd vdd FILL
XFILL_70_DFFSR_210 gnd vdd FILL
XFILL_70_DFFSR_221 gnd vdd FILL
XFILL_12_NAND3X1_103 gnd vdd FILL
XFILL_70_DFFSR_232 gnd vdd FILL
XFILL_70_DFFSR_243 gnd vdd FILL
XFILL_12_NAND3X1_114 gnd vdd FILL
XFILL_70_DFFSR_254 gnd vdd FILL
XFILL_12_NAND3X1_125 gnd vdd FILL
XFILL_11_3_1 gnd vdd FILL
XFILL_70_DFFSR_265 gnd vdd FILL
XFILL_24_NOR3X1_20 gnd vdd FILL
XFILL_24_NOR3X1_31 gnd vdd FILL
XFILL_24_NOR3X1_42 gnd vdd FILL
XFILL_74_DFFSR_220 gnd vdd FILL
XFILL_74_DFFSR_231 gnd vdd FILL
XFILL_74_DFFSR_242 gnd vdd FILL
XFILL_3_BUFX4_1 gnd vdd FILL
XFILL_74_DFFSR_253 gnd vdd FILL
XFILL_74_DFFSR_264 gnd vdd FILL
XFILL_74_DFFSR_275 gnd vdd FILL
XFILL_28_DFFSR_9 gnd vdd FILL
XFILL_28_NOR3X1_30 gnd vdd FILL
XFILL_28_NOR3X1_41 gnd vdd FILL
XFILL_13_MUX2X1_103 gnd vdd FILL
XFILL_5_CLKBUF1_40 gnd vdd FILL
XFILL_28_NOR3X1_52 gnd vdd FILL
XOAI22X1_1 INVX1_72/Y OAI22X1_1/B INVX1_76/Y OAI22X1_1/D gnd OAI22X1_1/Y vdd OAI22X1
XFILL_13_MUX2X1_114 gnd vdd FILL
XFILL_13_MUX2X1_125 gnd vdd FILL
XFILL_78_DFFSR_230 gnd vdd FILL
XFILL_7_OAI22X1_9 gnd vdd FILL
XFILL_3_NAND3X1_108 gnd vdd FILL
XFILL_13_MUX2X1_136 gnd vdd FILL
XFILL_78_DFFSR_241 gnd vdd FILL
XFILL_13_MUX2X1_147 gnd vdd FILL
XFILL_13_MUX2X1_158 gnd vdd FILL
XFILL_78_DFFSR_252 gnd vdd FILL
XFILL_3_NAND3X1_119 gnd vdd FILL
XFILL_0_AOI21X1_70 gnd vdd FILL
XFILL_78_DFFSR_263 gnd vdd FILL
XFILL_78_DFFSR_274 gnd vdd FILL
XFILL_33_CLKBUF1_4 gnd vdd FILL
XFILL_13_MUX2X1_169 gnd vdd FILL
XFILL_0_AOI21X1_81 gnd vdd FILL
XFILL_10_OAI22X1_50 gnd vdd FILL
XFILL_14_OAI21X1_30 gnd vdd FILL
XFILL_14_OAI21X1_41 gnd vdd FILL
XFILL_2_INVX1_5 gnd vdd FILL
XFILL_3_NOR2X1_180 gnd vdd FILL
XFILL_3_NOR2X1_191 gnd vdd FILL
XFILL_56_DFFSR_209 gnd vdd FILL
XFILL_19_4_1 gnd vdd FILL
XFILL_62_7_2 gnd vdd FILL
XFILL_83_DFFSR_109 gnd vdd FILL
XFILL_61_2_1 gnd vdd FILL
XFILL_21_5 gnd vdd FILL
XFILL_20_MUX2X1_160 gnd vdd FILL
XFILL_20_MUX2X1_171 gnd vdd FILL
XFILL_3_MUX2X1_120 gnd vdd FILL
XFILL_87_DFFSR_108 gnd vdd FILL
XFILL_20_MUX2X1_182 gnd vdd FILL
XFILL_3_INVX4_1 gnd vdd FILL
XFILL_14_4 gnd vdd FILL
XFILL_20_MUX2X1_193 gnd vdd FILL
XFILL_87_DFFSR_119 gnd vdd FILL
XFILL_3_MUX2X1_131 gnd vdd FILL
XFILL_14_BUFX4_13 gnd vdd FILL
XFILL_3_MUX2X1_142 gnd vdd FILL
XFILL_3_MUX2X1_153 gnd vdd FILL
XFILL_14_BUFX4_24 gnd vdd FILL
XFILL_3_MUX2X1_164 gnd vdd FILL
XFILL_14_BUFX4_35 gnd vdd FILL
XFILL_3_MUX2X1_175 gnd vdd FILL
XFILL_14_BUFX4_46 gnd vdd FILL
XFILL_14_BUFX4_57 gnd vdd FILL
XFILL_3_MUX2X1_186 gnd vdd FILL
XDFFSR_203 NOR2X1_28/A DFFSR_39/CLK DFFSR_45/R vdd DFFSR_203/D gnd vdd DFFSR
XFILL_14_BUFX4_68 gnd vdd FILL
XDFFSR_214 INVX1_81/A DFFSR_57/CLK DFFSR_90/R vdd MUX2X1_67/Y gnd vdd DFFSR
XDFFSR_225 INVX1_74/A DFFSR_47/CLK DFFSR_6/R vdd MUX2X1_61/Y gnd vdd DFFSR
XFILL_14_BUFX4_79 gnd vdd FILL
XDFFSR_236 INVX1_59/A CLKBUF1_5/Y BUFX4_23/Y vdd MUX2X1_45/Y gnd vdd DFFSR
XDFFSR_247 INVX1_52/A DFFSR_39/CLK DFFSR_45/R vdd MUX2X1_39/Y gnd vdd DFFSR
XDFFSR_258 NOR2X1_15/A DFFSR_6/CLK BUFX4_54/Y vdd DFFSR_258/D gnd vdd DFFSR
XFILL_41_DFFSR_220 gnd vdd FILL
XDFFSR_269 INVX1_38/A DFFSR_8/CLK DFFSR_9/R vdd MUX2X1_25/Y gnd vdd DFFSR
XFILL_41_DFFSR_231 gnd vdd FILL
XFILL_41_DFFSR_242 gnd vdd FILL
XFILL_41_DFFSR_253 gnd vdd FILL
XFILL_41_DFFSR_264 gnd vdd FILL
XFILL_41_DFFSR_275 gnd vdd FILL
XFILL_0_NOR2X1_90 gnd vdd FILL
XFILL_45_DFFSR_230 gnd vdd FILL
XFILL_45_DFFSR_241 gnd vdd FILL
XFILL_45_DFFSR_252 gnd vdd FILL
XFILL_45_DFFSR_263 gnd vdd FILL
XFILL_45_DFFSR_274 gnd vdd FILL
XFILL_72_DFFSR_130 gnd vdd FILL
XFILL_72_DFFSR_141 gnd vdd FILL
XFILL_9_AND2X2_6 gnd vdd FILL
XFILL_72_DFFSR_152 gnd vdd FILL
XFILL_49_DFFSR_240 gnd vdd FILL
XFILL_49_DFFSR_251 gnd vdd FILL
XFILL_49_DFFSR_262 gnd vdd FILL
XFILL_72_DFFSR_163 gnd vdd FILL
XFILL_72_DFFSR_174 gnd vdd FILL
XFILL_49_DFFSR_273 gnd vdd FILL
XFILL_72_DFFSR_185 gnd vdd FILL
XFILL_72_DFFSR_196 gnd vdd FILL
XFILL_23_DFFSR_209 gnd vdd FILL
XFILL_6_NAND3X1_12 gnd vdd FILL
XFILL_6_NAND3X1_23 gnd vdd FILL
XFILL_76_DFFSR_140 gnd vdd FILL
XFILL_6_NAND3X1_34 gnd vdd FILL
XFILL_53_7_2 gnd vdd FILL
XFILL_76_DFFSR_151 gnd vdd FILL
XFILL_6_NAND3X1_45 gnd vdd FILL
XFILL_76_DFFSR_162 gnd vdd FILL
XFILL_6_NAND3X1_56 gnd vdd FILL
XFILL_45_DFFSR_3 gnd vdd FILL
XFILL_52_2_1 gnd vdd FILL
XFILL_76_DFFSR_173 gnd vdd FILL
XFILL_6_NAND3X1_67 gnd vdd FILL
XFILL_6_BUFX4_12 gnd vdd FILL
XFILL_76_DFFSR_184 gnd vdd FILL
XFILL_6_NAND3X1_78 gnd vdd FILL
XFILL_6_BUFX4_23 gnd vdd FILL
XFILL_6_NAND3X1_89 gnd vdd FILL
XFILL_76_DFFSR_195 gnd vdd FILL
XFILL_50_DFFSR_109 gnd vdd FILL
XFILL_27_DFFSR_208 gnd vdd FILL
XFILL_6_BUFX4_34 gnd vdd FILL
XFILL_6_BUFX4_45 gnd vdd FILL
XFILL_27_DFFSR_219 gnd vdd FILL
XFILL_6_BUFX4_56 gnd vdd FILL
XFILL_66_10 gnd vdd FILL
XFILL_6_BUFX4_67 gnd vdd FILL
XFILL_6_BUFX4_78 gnd vdd FILL
XFILL_6_BUFX4_89 gnd vdd FILL
XFILL_0_NAND2X1_1 gnd vdd FILL
XFILL_54_DFFSR_108 gnd vdd FILL
XFILL_8_BUFX2_8 gnd vdd FILL
XFILL_54_DFFSR_119 gnd vdd FILL
XFILL_13_AOI21X1_19 gnd vdd FILL
XFILL_58_DFFSR_107 gnd vdd FILL
XFILL_58_DFFSR_118 gnd vdd FILL
XFILL_58_DFFSR_129 gnd vdd FILL
XFILL_67_DFFSR_7 gnd vdd FILL
XFILL_50_DFFSR_19 gnd vdd FILL
XFILL_12_DFFSR_230 gnd vdd FILL
XFILL_12_DFFSR_241 gnd vdd FILL
XFILL_12_DFFSR_252 gnd vdd FILL
XFILL_12_DFFSR_263 gnd vdd FILL
XFILL_12_DFFSR_274 gnd vdd FILL
XFILL_25_CLKBUF1_13 gnd vdd FILL
XFILL_25_CLKBUF1_24 gnd vdd FILL
XFILL_0_AOI21X1_6 gnd vdd FILL
XFILL_25_CLKBUF1_35 gnd vdd FILL
XFILL_10_BUFX4_50 gnd vdd FILL
XFILL_10_BUFX4_61 gnd vdd FILL
XFILL_16_DFFSR_240 gnd vdd FILL
XFILL_7_BUFX4_2 gnd vdd FILL
XFILL_16_DFFSR_251 gnd vdd FILL
XFILL_16_DFFSR_262 gnd vdd FILL
XFILL_10_BUFX4_72 gnd vdd FILL
XFILL_10_BUFX4_83 gnd vdd FILL
XFILL_9_DFFSR_109 gnd vdd FILL
XFILL_16_DFFSR_273 gnd vdd FILL
XFILL_8_CLKBUF1_17 gnd vdd FILL
XFILL_8_CLKBUF1_28 gnd vdd FILL
XFILL_10_BUFX4_94 gnd vdd FILL
XFILL_13_MUX2X1_18 gnd vdd FILL
XFILL_44_7_2 gnd vdd FILL
XFILL_13_MUX2X1_29 gnd vdd FILL
XFILL_8_CLKBUF1_39 gnd vdd FILL
XFILL_3_AOI21X1_14 gnd vdd FILL
XFILL_4_AOI21X1_5 gnd vdd FILL
XFILL_43_2_1 gnd vdd FILL
XFILL_3_AOI21X1_25 gnd vdd FILL
XFILL_43_DFFSR_140 gnd vdd FILL
XFILL_43_DFFSR_151 gnd vdd FILL
XFILL_3_AOI21X1_36 gnd vdd FILL
XFILL_3_AOI21X1_47 gnd vdd FILL
XFILL_43_DFFSR_162 gnd vdd FILL
XFILL_3_AOI21X1_58 gnd vdd FILL
XFILL_3_AOI21X1_69 gnd vdd FILL
XOAI21X1_17 INVX1_189/Y OAI21X1_7/B OAI21X1_17/C gnd NOR2X1_78/A vdd OAI21X1
XFILL_43_DFFSR_173 gnd vdd FILL
XFILL_13_OAI22X1_16 gnd vdd FILL
XFILL_43_DFFSR_184 gnd vdd FILL
XOAI21X1_28 INVX1_158/Y OAI21X1_3/B OAI21X1_28/C gnd OAI21X1_28/Y vdd OAI21X1
XFILL_13_OAI22X1_27 gnd vdd FILL
XFILL_43_DFFSR_195 gnd vdd FILL
XOAI21X1_39 INVX2_5/A OAI21X1_39/B OAI21X1_48/A gnd OAI21X1_39/Y vdd OAI21X1
XFILL_13_OAI22X1_38 gnd vdd FILL
XFILL_17_MUX2X1_17 gnd vdd FILL
XFILL_6_NOR2X1_102 gnd vdd FILL
XFILL_17_MUX2X1_28 gnd vdd FILL
XFILL_13_OAI22X1_49 gnd vdd FILL
XFILL_6_NOR2X1_113 gnd vdd FILL
XFILL_17_MUX2X1_39 gnd vdd FILL
XFILL_8_AOI21X1_4 gnd vdd FILL
XFILL_6_NOR2X1_124 gnd vdd FILL
XFILL_2_DFFSR_19 gnd vdd FILL
XFILL_47_DFFSR_150 gnd vdd FILL
XFILL_6_NOR2X1_135 gnd vdd FILL
XFILL_47_DFFSR_161 gnd vdd FILL
XFILL_6_NOR2X1_146 gnd vdd FILL
XFILL_13_NAND3X1_104 gnd vdd FILL
XFILL_6_NOR2X1_157 gnd vdd FILL
XFILL_13_NAND3X1_115 gnd vdd FILL
XFILL_47_DFFSR_172 gnd vdd FILL
XFILL_6_INVX1_6 gnd vdd FILL
XFILL_47_DFFSR_183 gnd vdd FILL
XFILL_13_NAND3X1_126 gnd vdd FILL
XFILL_6_NOR2X1_168 gnd vdd FILL
XFILL_6_NOR2X1_179 gnd vdd FILL
XFILL_47_DFFSR_194 gnd vdd FILL
XFILL_21_DFFSR_108 gnd vdd FILL
XFILL_12_NAND3X1_70 gnd vdd FILL
XFILL_12_NAND3X1_81 gnd vdd FILL
XFILL_21_DFFSR_119 gnd vdd FILL
XFILL_4_INVX1_40 gnd vdd FILL
XFILL_4_INVX1_51 gnd vdd FILL
XFILL_12_NAND3X1_92 gnd vdd FILL
XFILL_4_INVX1_62 gnd vdd FILL
XFILL_13_AOI22X1_1 gnd vdd FILL
XFILL_4_INVX1_73 gnd vdd FILL
XFILL_4_INVX1_84 gnd vdd FILL
XFILL_4_INVX1_95 gnd vdd FILL
XFILL_25_DFFSR_107 gnd vdd FILL
XFILL_23_MUX2X1_104 gnd vdd FILL
XFILL_11_MUX2X1_5 gnd vdd FILL
XFILL_25_DFFSR_118 gnd vdd FILL
XFILL_25_DFFSR_129 gnd vdd FILL
XFILL_23_MUX2X1_115 gnd vdd FILL
XFILL_23_MUX2X1_126 gnd vdd FILL
XFILL_23_MUX2X1_137 gnd vdd FILL
XFILL_4_NAND3X1_109 gnd vdd FILL
XFILL_23_MUX2X1_148 gnd vdd FILL
XFILL_23_MUX2X1_159 gnd vdd FILL
XFILL_29_DFFSR_106 gnd vdd FILL
XFILL_6_MUX2X1_108 gnd vdd FILL
XFILL_6_MUX2X1_119 gnd vdd FILL
XFILL_2_BUFX4_60 gnd vdd FILL
XFILL_29_DFFSR_117 gnd vdd FILL
XFILL_19_DFFSR_20 gnd vdd FILL
XFILL_2_BUFX4_71 gnd vdd FILL
XFILL_19_DFFSR_31 gnd vdd FILL
XFILL_29_DFFSR_128 gnd vdd FILL
XFILL_19_DFFSR_42 gnd vdd FILL
XFILL_29_DFFSR_139 gnd vdd FILL
XFILL_19_DFFSR_53 gnd vdd FILL
XFILL_3_OAI22X1_11 gnd vdd FILL
XFILL_2_BUFX4_82 gnd vdd FILL
XFILL_2_BUFX4_93 gnd vdd FILL
XFILL_3_OAI22X1_22 gnd vdd FILL
XFILL_19_DFFSR_64 gnd vdd FILL
XFILL_19_DFFSR_75 gnd vdd FILL
XFILL_3_OAI22X1_33 gnd vdd FILL
XFILL_3_OAI22X1_44 gnd vdd FILL
XFILL_19_DFFSR_86 gnd vdd FILL
XFILL_21_NOR3X1_19 gnd vdd FILL
XFILL_19_DFFSR_97 gnd vdd FILL
XFILL_7_OAI21X1_13 gnd vdd FILL
XFILL_7_OAI21X1_24 gnd vdd FILL
XFILL_71_DFFSR_208 gnd vdd FILL
XFILL_59_DFFSR_30 gnd vdd FILL
XFILL_7_OAI21X1_35 gnd vdd FILL
XFILL_71_DFFSR_219 gnd vdd FILL
XFILL_59_DFFSR_41 gnd vdd FILL
XFILL_7_OAI21X1_46 gnd vdd FILL
XFILL_59_DFFSR_52 gnd vdd FILL
XFILL_59_DFFSR_63 gnd vdd FILL
XFILL_20_MUX2X1_3 gnd vdd FILL
XFILL_35_7_2 gnd vdd FILL
XFILL_59_DFFSR_74 gnd vdd FILL
XFILL_25_NOR3X1_18 gnd vdd FILL
XFILL_59_DFFSR_85 gnd vdd FILL
XFILL_34_2_1 gnd vdd FILL
XFILL_59_DFFSR_96 gnd vdd FILL
XFILL_25_NOR3X1_29 gnd vdd FILL
XFILL_75_DFFSR_207 gnd vdd FILL
XFILL_0_NOR2X1_202 gnd vdd FILL
XFILL_4_NOR2X1_6 gnd vdd FILL
XFILL_84_DFFSR_1 gnd vdd FILL
XFILL_75_DFFSR_218 gnd vdd FILL
XFILL_10_DFFSR_140 gnd vdd FILL
XFILL_10_DFFSR_151 gnd vdd FILL
XFILL_75_DFFSR_229 gnd vdd FILL
XFILL_10_DFFSR_162 gnd vdd FILL
XFILL_28_DFFSR_40 gnd vdd FILL
XFILL_29_NOR3X1_17 gnd vdd FILL
XFILL_10_DFFSR_173 gnd vdd FILL
XFILL_12_1 gnd vdd FILL
XFILL_10_DFFSR_184 gnd vdd FILL
XFILL_28_DFFSR_51 gnd vdd FILL
XFILL_29_NOR3X1_28 gnd vdd FILL
XFILL_28_DFFSR_62 gnd vdd FILL
XFILL_29_NOR3X1_39 gnd vdd FILL
XFILL_10_DFFSR_195 gnd vdd FILL
XFILL_28_DFFSR_73 gnd vdd FILL
XFILL_79_DFFSR_206 gnd vdd FILL
XFILL_28_DFFSR_84 gnd vdd FILL
XFILL_14_CLKBUF1_20 gnd vdd FILL
XFILL_79_DFFSR_217 gnd vdd FILL
XFILL_14_CLKBUF1_31 gnd vdd FILL
XFILL_28_DFFSR_95 gnd vdd FILL
XFILL_14_CLKBUF1_42 gnd vdd FILL
XFILL_79_DFFSR_228 gnd vdd FILL
XFILL_14_DFFSR_150 gnd vdd FILL
XFILL_14_DFFSR_161 gnd vdd FILL
XFILL_79_DFFSR_239 gnd vdd FILL
XFILL_14_DFFSR_172 gnd vdd FILL
XFILL_3_CLKBUF1_4 gnd vdd FILL
XFILL_3_MUX2X1_4 gnd vdd FILL
XFILL_14_DFFSR_183 gnd vdd FILL
XFILL_68_DFFSR_50 gnd vdd FILL
XFILL_14_DFFSR_194 gnd vdd FILL
XFILL_68_DFFSR_61 gnd vdd FILL
XFILL_68_DFFSR_72 gnd vdd FILL
XFILL_68_DFFSR_83 gnd vdd FILL
XFILL_11_DFFSR_6 gnd vdd FILL
XFILL_68_DFFSR_94 gnd vdd FILL
XFILL_18_DFFSR_160 gnd vdd FILL
XFILL_49_DFFSR_4 gnd vdd FILL
XFILL_7_CLKBUF1_3 gnd vdd FILL
XFILL_18_DFFSR_171 gnd vdd FILL
XFILL_18_DFFSR_182 gnd vdd FILL
XFILL_18_DFFSR_193 gnd vdd FILL
XFILL_10_NOR3X1_40 gnd vdd FILL
XFILL_10_NOR3X1_51 gnd vdd FILL
XFILL_37_DFFSR_60 gnd vdd FILL
XFILL_37_DFFSR_71 gnd vdd FILL
XFILL_37_DFFSR_82 gnd vdd FILL
XFILL_60_DFFSR_240 gnd vdd FILL
XFILL_37_DFFSR_93 gnd vdd FILL
XFILL_60_DFFSR_251 gnd vdd FILL
XFILL_60_DFFSR_262 gnd vdd FILL
XFILL_60_DFFSR_273 gnd vdd FILL
XFILL_14_NOR3X1_50 gnd vdd FILL
XFILL_77_DFFSR_70 gnd vdd FILL
XFILL_77_DFFSR_81 gnd vdd FILL
XFILL_77_DFFSR_92 gnd vdd FILL
XFILL_64_DFFSR_250 gnd vdd FILL
XFILL_64_DFFSR_261 gnd vdd FILL
XFILL_64_DFFSR_272 gnd vdd FILL
XFILL_12_MUX2X1_100 gnd vdd FILL
XFILL_26_7_2 gnd vdd FILL
XFILL_12_MUX2X1_111 gnd vdd FILL
XFILL_1_7_2 gnd vdd FILL
XFILL_12_MUX2X1_122 gnd vdd FILL
XFILL_0_OAI21X1_9 gnd vdd FILL
XFILL_25_2_1 gnd vdd FILL
XFILL_0_2_1 gnd vdd FILL
XFILL_12_MUX2X1_133 gnd vdd FILL
XFILL_12_MUX2X1_144 gnd vdd FILL
XFILL_12_MUX2X1_155 gnd vdd FILL
XFILL_68_DFFSR_260 gnd vdd FILL
XFILL_68_DFFSR_271 gnd vdd FILL
XFILL_23_CLKBUF1_1 gnd vdd FILL
XFILL_12_MUX2X1_166 gnd vdd FILL
XFILL_12_MUX2X1_177 gnd vdd FILL
XFILL_46_DFFSR_80 gnd vdd FILL
XFILL_12_MUX2X1_188 gnd vdd FILL
XFILL_1_NOR2X1_11 gnd vdd FILL
XFILL_42_DFFSR_207 gnd vdd FILL
XFILL_46_DFFSR_91 gnd vdd FILL
XFILL_42_DFFSR_218 gnd vdd FILL
XFILL_1_NOR2X1_22 gnd vdd FILL
XFILL_4_OAI21X1_8 gnd vdd FILL
XFILL_1_NOR2X1_33 gnd vdd FILL
XFILL_1_NOR2X1_44 gnd vdd FILL
XFILL_42_DFFSR_229 gnd vdd FILL
XFILL_1_NOR2X1_55 gnd vdd FILL
XFILL_1_NOR2X1_66 gnd vdd FILL
XFILL_1_NOR2X1_77 gnd vdd FILL
XFILL_1_NOR2X1_88 gnd vdd FILL
XFILL_1_NOR2X1_99 gnd vdd FILL
XFILL_5_NOR2X1_10 gnd vdd FILL
XFILL_46_DFFSR_206 gnd vdd FILL
XFILL_86_DFFSR_90 gnd vdd FILL
XFILL_5_NOR2X1_21 gnd vdd FILL
XFILL_46_DFFSR_217 gnd vdd FILL
XFILL_8_OAI21X1_7 gnd vdd FILL
XFILL_46_DFFSR_228 gnd vdd FILL
XFILL_5_NOR2X1_32 gnd vdd FILL
XFILL_5_NOR2X1_43 gnd vdd FILL
XFILL_5_NOR2X1_54 gnd vdd FILL
XFILL_46_DFFSR_239 gnd vdd FILL
XFILL_15_DFFSR_90 gnd vdd FILL
XFILL_5_NOR2X1_65 gnd vdd FILL
XFILL_5_NOR2X1_76 gnd vdd FILL
XFILL_5_NOR2X1_87 gnd vdd FILL
XFILL_73_DFFSR_106 gnd vdd FILL
XFILL_5_NOR2X1_98 gnd vdd FILL
XFILL_9_NOR2X1_20 gnd vdd FILL
XFILL_73_DFFSR_117 gnd vdd FILL
XFILL_9_NOR2X1_31 gnd vdd FILL
XFILL_73_DFFSR_128 gnd vdd FILL
XFILL_9_NOR2X1_42 gnd vdd FILL
XFILL_73_DFFSR_139 gnd vdd FILL
XFILL_9_NOR2X1_53 gnd vdd FILL
XFILL_13_OAI22X1_4 gnd vdd FILL
XFILL_9_NOR2X1_64 gnd vdd FILL
XFILL_9_NOR2X1_75 gnd vdd FILL
XFILL_9_NOR2X1_86 gnd vdd FILL
XFILL_77_DFFSR_105 gnd vdd FILL
XFILL_8_3_1 gnd vdd FILL
XFILL_9_NOR2X1_97 gnd vdd FILL
XFILL_77_DFFSR_116 gnd vdd FILL
XFILL_77_DFFSR_127 gnd vdd FILL
XFILL_77_DFFSR_138 gnd vdd FILL
XFILL_2_MUX2X1_150 gnd vdd FILL
XFILL_2_MUX2X1_161 gnd vdd FILL
XFILL_77_DFFSR_149 gnd vdd FILL
XFILL_17_OAI22X1_3 gnd vdd FILL
XFILL_15_NAND3X1_14 gnd vdd FILL
XFILL_15_NAND3X1_25 gnd vdd FILL
XFILL_2_MUX2X1_172 gnd vdd FILL
XFILL_2_MUX2X1_183 gnd vdd FILL
XFILL_15_NAND3X1_36 gnd vdd FILL
XFILL_2_MUX2X1_194 gnd vdd FILL
XFILL_15_NAND3X1_47 gnd vdd FILL
XFILL_15_NAND3X1_58 gnd vdd FILL
XFILL_15_NAND3X1_69 gnd vdd FILL
XFILL_35_CLKBUF1_14 gnd vdd FILL
XFILL_35_CLKBUF1_25 gnd vdd FILL
XFILL_35_CLKBUF1_36 gnd vdd FILL
XFILL_17_7_2 gnd vdd FILL
XFILL_31_DFFSR_250 gnd vdd FILL
XFILL_31_DFFSR_261 gnd vdd FILL
XFILL_31_DFFSR_272 gnd vdd FILL
XFILL_16_2_1 gnd vdd FILL
XFILL_11_BUFX4_17 gnd vdd FILL
XFILL_11_BUFX4_28 gnd vdd FILL
XFILL_35_DFFSR_260 gnd vdd FILL
XFILL_35_DFFSR_271 gnd vdd FILL
XFILL_11_BUFX4_39 gnd vdd FILL
XFILL_5_NAND2X1_9 gnd vdd FILL
XFILL_1_MUX2X1_40 gnd vdd FILL
XFILL_1_MUX2X1_51 gnd vdd FILL
XFILL_1_MUX2X1_62 gnd vdd FILL
XFILL_1_MUX2X1_73 gnd vdd FILL
XFILL_62_DFFSR_160 gnd vdd FILL
XFILL_1_MUX2X1_84 gnd vdd FILL
XFILL_14_NAND3X1_105 gnd vdd FILL
XFILL_1_MUX2X1_95 gnd vdd FILL
XFILL_14_NAND3X1_116 gnd vdd FILL
XFILL_39_DFFSR_270 gnd vdd FILL
XFILL_14_NAND3X1_127 gnd vdd FILL
XFILL_62_DFFSR_171 gnd vdd FILL
XFILL_62_DFFSR_182 gnd vdd FILL
XFILL_62_DFFSR_193 gnd vdd FILL
XFILL_9_NAND2X1_8 gnd vdd FILL
XFILL_13_DFFSR_206 gnd vdd FILL
XFILL_13_DFFSR_217 gnd vdd FILL
XFILL_10_NAND3X1_6 gnd vdd FILL
XFILL_5_MUX2X1_50 gnd vdd FILL
XFILL_5_NAND3X1_20 gnd vdd FILL
XFILL_5_MUX2X1_61 gnd vdd FILL
XFILL_13_DFFSR_228 gnd vdd FILL
XFILL_5_NAND3X1_31 gnd vdd FILL
XFILL_5_MUX2X1_72 gnd vdd FILL
XFILL_13_DFFSR_239 gnd vdd FILL
XFILL_5_NAND3X1_42 gnd vdd FILL
XFILL_5_MUX2X1_83 gnd vdd FILL
XFILL_5_NAND3X1_53 gnd vdd FILL
XFILL_50_DFFSR_4 gnd vdd FILL
XFILL_66_DFFSR_170 gnd vdd FILL
XFILL_5_MUX2X1_94 gnd vdd FILL
XFILL_9_NAND2X1_11 gnd vdd FILL
XFILL_5_NAND3X1_64 gnd vdd FILL
XFILL_9_NAND2X1_22 gnd vdd FILL
XFILL_5_NAND3X1_75 gnd vdd FILL
XFILL_66_DFFSR_181 gnd vdd FILL
XFILL_9_NAND2X1_33 gnd vdd FILL
XFILL_5_NAND3X1_86 gnd vdd FILL
XFILL_66_DFFSR_192 gnd vdd FILL
XFILL_40_DFFSR_106 gnd vdd FILL
XFILL_17_DFFSR_205 gnd vdd FILL
XFILL_9_NAND2X1_44 gnd vdd FILL
XFILL_5_NAND3X1_97 gnd vdd FILL
XFILL_9_NAND2X1_55 gnd vdd FILL
XFILL_17_DFFSR_216 gnd vdd FILL
XFILL_40_DFFSR_117 gnd vdd FILL
XFILL_14_NAND3X1_5 gnd vdd FILL
XFILL_9_NAND2X1_66 gnd vdd FILL
XFILL_17_DFFSR_227 gnd vdd FILL
XFILL_9_MUX2X1_60 gnd vdd FILL
XFILL_40_DFFSR_128 gnd vdd FILL
XFILL_9_MUX2X1_71 gnd vdd FILL
XFILL_9_NAND2X1_77 gnd vdd FILL
XFILL_40_DFFSR_139 gnd vdd FILL
XFILL_17_DFFSR_238 gnd vdd FILL
XFILL_5_INVX1_18 gnd vdd FILL
XFILL_9_MUX2X1_82 gnd vdd FILL
XFILL_9_NAND2X1_88 gnd vdd FILL
XFILL_22_15 gnd vdd FILL
XCLKBUF1_18 BUFX4_10/Y gnd DFFSR_93/CLK vdd CLKBUF1
XFILL_5_INVX1_29 gnd vdd FILL
XFILL_17_DFFSR_249 gnd vdd FILL
XFILL_9_MUX2X1_93 gnd vdd FILL
XCLKBUF1_29 BUFX4_84/Y gnd DFFSR_72/CLK vdd CLKBUF1
XFILL_44_DFFSR_105 gnd vdd FILL
XFILL_67_2 gnd vdd FILL
XFILL_17_CLKBUF1_19 gnd vdd FILL
XFILL_44_DFFSR_116 gnd vdd FILL
XFILL_44_DFFSR_127 gnd vdd FILL
XFILL_44_DFFSR_138 gnd vdd FILL
XBUFX4_50 BUFX4_51/Y gnd BUFX4_50/Y vdd BUFX4
XFILL_66_1_1 gnd vdd FILL
XFILL_44_DFFSR_149 gnd vdd FILL
XBUFX4_61 INVX8_1/Y gnd MUX2X1_9/A vdd BUFX4
XFILL_12_AOI21X1_16 gnd vdd FILL
XFILL_12_AOI21X1_27 gnd vdd FILL
XBUFX4_72 INVX8_2/Y gnd BUFX4_72/Y vdd BUFX4
XBUFX4_83 INVX8_4/Y gnd BUFX4_83/Y vdd BUFX4
XFILL_12_AOI21X1_38 gnd vdd FILL
XFILL_12_AOI21X1_49 gnd vdd FILL
XFILL_2_DFFSR_9 gnd vdd FILL
XBUFX4_94 INVX8_3/Y gnd MUX2X1_7/B vdd BUFX4
XFILL_48_DFFSR_104 gnd vdd FILL
XFILL_48_DFFSR_115 gnd vdd FILL
XFILL_15_DFFSR_7 gnd vdd FILL
XFILL_3_BUFX4_16 gnd vdd FILL
XFILL_48_DFFSR_126 gnd vdd FILL
XFILL_48_DFFSR_137 gnd vdd FILL
XFILL_3_BUFX4_27 gnd vdd FILL
XFILL_72_DFFSR_8 gnd vdd FILL
XFILL_48_DFFSR_148 gnd vdd FILL
XFILL_3_BUFX4_38 gnd vdd FILL
XFILL_48_DFFSR_159 gnd vdd FILL
XFILL_3_BUFX4_49 gnd vdd FILL
XFILL_21_MUX2X1_70 gnd vdd FILL
XFILL_21_MUX2X1_81 gnd vdd FILL
XFILL_21_MUX2X1_92 gnd vdd FILL
XFILL_50_5_2 gnd vdd FILL
XFILL_24_CLKBUF1_10 gnd vdd FILL
XFILL_24_CLKBUF1_21 gnd vdd FILL
XFILL_24_CLKBUF1_32 gnd vdd FILL
XFILL_0_NAND3X1_106 gnd vdd FILL
XFILL_18_AOI22X1_9 gnd vdd FILL
XFILL_0_NAND3X1_117 gnd vdd FILL
XFILL_0_NAND3X1_128 gnd vdd FILL
XFILL_7_CLKBUF1_14 gnd vdd FILL
XFILL_7_CLKBUF1_25 gnd vdd FILL
XFILL_10_AND2X2_4 gnd vdd FILL
XFILL_7_CLKBUF1_36 gnd vdd FILL
XFILL_29_DFFSR_18 gnd vdd FILL
XFILL_2_AOI21X1_11 gnd vdd FILL
XFILL_29_DFFSR_29 gnd vdd FILL
XFILL_2_AOI21X1_22 gnd vdd FILL
XFILL_2_AOI21X1_33 gnd vdd FILL
XFILL_2_AOI21X1_44 gnd vdd FILL
XFILL_2_AOI21X1_55 gnd vdd FILL
XFILL_12_OAI22X1_13 gnd vdd FILL
XFILL_33_DFFSR_170 gnd vdd FILL
XFILL_2_AOI21X1_66 gnd vdd FILL
XFILL_2_AOI21X1_77 gnd vdd FILL
XFILL_12_OAI22X1_24 gnd vdd FILL
XFILL_33_DFFSR_181 gnd vdd FILL
XFILL_12_OAI22X1_35 gnd vdd FILL
XFILL_69_DFFSR_17 gnd vdd FILL
XFILL_33_DFFSR_192 gnd vdd FILL
XFILL_12_OAI22X1_46 gnd vdd FILL
XFILL_69_DFFSR_28 gnd vdd FILL
XFILL_5_NOR2X1_110 gnd vdd FILL
XFILL_69_DFFSR_39 gnd vdd FILL
XFILL_5_NOR2X1_121 gnd vdd FILL
XFILL_5_NOR2X1_132 gnd vdd FILL
XFILL_5_NOR2X1_143 gnd vdd FILL
XFILL_58_6_2 gnd vdd FILL
XFILL_5_NOR2X1_154 gnd vdd FILL
XFILL_5_NOR2X1_165 gnd vdd FILL
XFILL_37_DFFSR_180 gnd vdd FILL
XFILL_57_1_1 gnd vdd FILL
XFILL_11_DFFSR_105 gnd vdd FILL
XFILL_5_NOR2X1_176 gnd vdd FILL
XFILL_37_DFFSR_191 gnd vdd FILL
XFILL_5_NOR2X1_187 gnd vdd FILL
XFILL_5_NOR2X1_198 gnd vdd FILL
XFILL_11_DFFSR_116 gnd vdd FILL
XFILL_11_DFFSR_127 gnd vdd FILL
XFILL_11_DFFSR_138 gnd vdd FILL
XFILL_11_DFFSR_149 gnd vdd FILL
XFILL_38_DFFSR_16 gnd vdd FILL
XFILL_38_DFFSR_27 gnd vdd FILL
XFILL_38_DFFSR_38 gnd vdd FILL
XFILL_38_DFFSR_49 gnd vdd FILL
XFILL_15_DFFSR_104 gnd vdd FILL
XFILL_15_DFFSR_115 gnd vdd FILL
XFILL_22_MUX2X1_101 gnd vdd FILL
XFILL_22_MUX2X1_112 gnd vdd FILL
XFILL_15_DFFSR_126 gnd vdd FILL
XFILL_15_DFFSR_137 gnd vdd FILL
XFILL_22_MUX2X1_123 gnd vdd FILL
XFILL_15_DFFSR_148 gnd vdd FILL
XFILL_78_DFFSR_15 gnd vdd FILL
XFILL_78_DFFSR_26 gnd vdd FILL
XFILL_15_DFFSR_159 gnd vdd FILL
XFILL_22_MUX2X1_134 gnd vdd FILL
XFILL_22_MUX2X1_145 gnd vdd FILL
XFILL_78_DFFSR_37 gnd vdd FILL
XFILL_22_MUX2X1_156 gnd vdd FILL
XFILL_41_5_2 gnd vdd FILL
XFILL_78_DFFSR_48 gnd vdd FILL
XFILL_22_MUX2X1_167 gnd vdd FILL
XFILL_83_DFFSR_270 gnd vdd FILL
XFILL_40_0_1 gnd vdd FILL
XFILL_19_DFFSR_103 gnd vdd FILL
XFILL_5_MUX2X1_105 gnd vdd FILL
XFILL_78_DFFSR_59 gnd vdd FILL
XFILL_5_MUX2X1_116 gnd vdd FILL
XFILL_19_DFFSR_114 gnd vdd FILL
XFILL_22_MUX2X1_178 gnd vdd FILL
XFILL_22_MUX2X1_189 gnd vdd FILL
XFILL_5_MUX2X1_127 gnd vdd FILL
XFILL_1_INVX1_11 gnd vdd FILL
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XFILL_1_INVX1_22 gnd vdd FILL
XFILL_19_DFFSR_125 gnd vdd FILL
XFILL_19_DFFSR_136 gnd vdd FILL
XFILL_5_MUX2X1_138 gnd vdd FILL
XFILL_1_INVX1_33 gnd vdd FILL
XFILL_5_MUX2X1_149 gnd vdd FILL
XFILL_19_DFFSR_147 gnd vdd FILL
XFILL_19_DFFSR_158 gnd vdd FILL
XFILL_1_INVX1_44 gnd vdd FILL
XFILL_2_AND2X2_3 gnd vdd FILL
XFILL_2_OAI22X1_30 gnd vdd FILL
XFILL_1_INVX1_55 gnd vdd FILL
XFILL_19_DFFSR_169 gnd vdd FILL
XFILL_1_INVX1_66 gnd vdd FILL
XFILL_11_NOR3X1_16 gnd vdd FILL
XFILL_2_OAI22X1_41 gnd vdd FILL
XFILL_1_INVX1_77 gnd vdd FILL
XFILL_1_INVX1_88 gnd vdd FILL
XFILL_11_NOR3X1_27 gnd vdd FILL
XFILL_6_OAI21X1_10 gnd vdd FILL
XFILL_47_DFFSR_14 gnd vdd FILL
XFILL_47_DFFSR_25 gnd vdd FILL
XFILL_6_OAI21X1_21 gnd vdd FILL
XFILL_1_INVX1_99 gnd vdd FILL
XFILL_47_DFFSR_36 gnd vdd FILL
XFILL_11_NOR3X1_38 gnd vdd FILL
XFILL_11_NOR3X1_49 gnd vdd FILL
XFILL_61_DFFSR_205 gnd vdd FILL
XFILL_6_OAI21X1_32 gnd vdd FILL
XFILL_47_DFFSR_47 gnd vdd FILL
XFILL_47_DFFSR_58 gnd vdd FILL
XFILL_61_DFFSR_216 gnd vdd FILL
XFILL_6_OAI21X1_43 gnd vdd FILL
XFILL_61_DFFSR_227 gnd vdd FILL
XFILL_47_DFFSR_69 gnd vdd FILL
XFILL_61_DFFSR_238 gnd vdd FILL
XFILL_61_DFFSR_249 gnd vdd FILL
XFILL_87_DFFSR_13 gnd vdd FILL
XFILL_15_NOR3X1_15 gnd vdd FILL
XFILL_15_NOR3X1_26 gnd vdd FILL
XFILL_87_DFFSR_24 gnd vdd FILL
XFILL_32_DFFSR_1 gnd vdd FILL
XFILL_15_NOR3X1_37 gnd vdd FILL
XFILL_87_DFFSR_35 gnd vdd FILL
XFILL_87_DFFSR_46 gnd vdd FILL
XFILL_15_NOR3X1_48 gnd vdd FILL
XFILL_65_DFFSR_204 gnd vdd FILL
XFILL_16_DFFSR_13 gnd vdd FILL
XFILL_65_DFFSR_215 gnd vdd FILL
XFILL_87_DFFSR_57 gnd vdd FILL
XFILL_87_DFFSR_68 gnd vdd FILL
XFILL_65_DFFSR_226 gnd vdd FILL
XFILL_16_DFFSR_24 gnd vdd FILL
XFILL_16_DFFSR_35 gnd vdd FILL
XFILL_65_DFFSR_237 gnd vdd FILL
XFILL_87_DFFSR_79 gnd vdd FILL
XFILL_16_DFFSR_46 gnd vdd FILL
XFILL_65_DFFSR_248 gnd vdd FILL
XFILL_19_NOR3X1_14 gnd vdd FILL
XFILL_16_DFFSR_57 gnd vdd FILL
XFILL_65_DFFSR_259 gnd vdd FILL
XFILL_16_DFFSR_68 gnd vdd FILL
XFILL_19_NOR3X1_25 gnd vdd FILL
XFILL_19_NOR3X1_36 gnd vdd FILL
XFILL_19_NOR3X1_47 gnd vdd FILL
XFILL_16_DFFSR_79 gnd vdd FILL
XFILL_49_6_2 gnd vdd FILL
XFILL_69_DFFSR_203 gnd vdd FILL
XFILL_60_9 gnd vdd FILL
XFILL_56_DFFSR_12 gnd vdd FILL
XFILL_69_DFFSR_214 gnd vdd FILL
XFILL_56_DFFSR_23 gnd vdd FILL
XFILL_69_DFFSR_225 gnd vdd FILL
XFILL_48_1_1 gnd vdd FILL
XFILL_69_DFFSR_236 gnd vdd FILL
XFILL_56_DFFSR_34 gnd vdd FILL
XFILL_27_NOR3X1_9 gnd vdd FILL
XFILL_69_DFFSR_247 gnd vdd FILL
XFILL_56_DFFSR_45 gnd vdd FILL
XFILL_56_DFFSR_56 gnd vdd FILL
XFILL_69_DFFSR_258 gnd vdd FILL
XFILL_69_DFFSR_269 gnd vdd FILL
XFILL_56_DFFSR_67 gnd vdd FILL
XFILL_56_DFFSR_78 gnd vdd FILL
XFILL_56_DFFSR_89 gnd vdd FILL
XFILL_8_NAND3X1_19 gnd vdd FILL
XFILL_54_DFFSR_5 gnd vdd FILL
XFILL_25_DFFSR_11 gnd vdd FILL
XFILL_25_DFFSR_22 gnd vdd FILL
XFILL_28_CLKBUF1_9 gnd vdd FILL
XFILL_25_DFFSR_33 gnd vdd FILL
XFILL_6_NOR2X1_19 gnd vdd FILL
XFILL_25_DFFSR_44 gnd vdd FILL
XFILL_25_DFFSR_55 gnd vdd FILL
XFILL_32_5_2 gnd vdd FILL
XFILL_25_DFFSR_66 gnd vdd FILL
XFILL_11_NOR2X1_190 gnd vdd FILL
XFILL_25_DFFSR_77 gnd vdd FILL
XFILL_25_DFFSR_88 gnd vdd FILL
XFILL_31_0_1 gnd vdd FILL
XFILL_25_DFFSR_99 gnd vdd FILL
XFILL_65_DFFSR_10 gnd vdd FILL
XFILL_65_DFFSR_21 gnd vdd FILL
XFILL_50_DFFSR_270 gnd vdd FILL
XFILL_65_DFFSR_32 gnd vdd FILL
XFILL_65_DFFSR_43 gnd vdd FILL
XFILL_0_MUX2X1_8 gnd vdd FILL
XFILL_65_DFFSR_54 gnd vdd FILL
XFILL_65_DFFSR_65 gnd vdd FILL
XFILL_65_DFFSR_76 gnd vdd FILL
XFILL_65_DFFSR_87 gnd vdd FILL
XFILL_65_DFFSR_98 gnd vdd FILL
XFILL_15_NAND3X1_106 gnd vdd FILL
XFILL_15_NAND3X1_117 gnd vdd FILL
XFILL_15_NAND3X1_128 gnd vdd FILL
XFILL_8_DFFSR_12 gnd vdd FILL
XFILL_8_DFFSR_23 gnd vdd FILL
XFILL_19_DFFSR_8 gnd vdd FILL
XFILL_8_DFFSR_34 gnd vdd FILL
XFILL_76_DFFSR_9 gnd vdd FILL
XFILL_34_DFFSR_20 gnd vdd FILL
XFILL_8_DFFSR_45 gnd vdd FILL
XFILL_8_DFFSR_56 gnd vdd FILL
XFILL_34_DFFSR_31 gnd vdd FILL
XFILL_8_DFFSR_67 gnd vdd FILL
XFILL_34_DFFSR_42 gnd vdd FILL
XFILL_11_MUX2X1_130 gnd vdd FILL
XFILL_8_DFFSR_78 gnd vdd FILL
XFILL_11_MUX2X1_141 gnd vdd FILL
XFILL_34_DFFSR_53 gnd vdd FILL
XFILL_8_DFFSR_89 gnd vdd FILL
XFILL_11_MUX2X1_152 gnd vdd FILL
XFILL_11_MUX2X1_163 gnd vdd FILL
XFILL_34_DFFSR_64 gnd vdd FILL
XFILL_34_DFFSR_75 gnd vdd FILL
XFILL_81_DFFSR_180 gnd vdd FILL
XFILL_34_DFFSR_86 gnd vdd FILL
XFILL_11_MUX2X1_174 gnd vdd FILL
XFILL_11_MUX2X1_185 gnd vdd FILL
XFILL_81_DFFSR_191 gnd vdd FILL
XFILL_34_DFFSR_97 gnd vdd FILL
XFILL_32_DFFSR_204 gnd vdd FILL
XFILL_32_DFFSR_215 gnd vdd FILL
XFILL_74_DFFSR_30 gnd vdd FILL
XFILL_32_DFFSR_226 gnd vdd FILL
XFILL_74_DFFSR_41 gnd vdd FILL
XFILL_32_DFFSR_237 gnd vdd FILL
XFILL_74_DFFSR_52 gnd vdd FILL
XFILL_1_DFFSR_250 gnd vdd FILL
XFILL_74_DFFSR_63 gnd vdd FILL
XFILL_32_DFFSR_248 gnd vdd FILL
XFILL_1_DFFSR_261 gnd vdd FILL
XFILL_1_DFFSR_272 gnd vdd FILL
XFILL_32_DFFSR_259 gnd vdd FILL
XFILL_74_DFFSR_74 gnd vdd FILL
XFILL_74_DFFSR_85 gnd vdd FILL
XFILL_85_DFFSR_190 gnd vdd FILL
XFILL_39_1_1 gnd vdd FILL
XFILL_74_DFFSR_96 gnd vdd FILL
XFILL_36_DFFSR_203 gnd vdd FILL
XFILL_36_DFFSR_214 gnd vdd FILL
XFILL_36_DFFSR_225 gnd vdd FILL
XFILL_36_DFFSR_236 gnd vdd FILL
XFILL_36_DFFSR_247 gnd vdd FILL
XFILL_5_DFFSR_260 gnd vdd FILL
XFILL_5_DFFSR_271 gnd vdd FILL
XFILL_36_DFFSR_258 gnd vdd FILL
XFILL_36_DFFSR_269 gnd vdd FILL
XFILL_2_MUX2X1_16 gnd vdd FILL
XFILL_43_DFFSR_40 gnd vdd FILL
XFILL_14_NOR3X1_4 gnd vdd FILL
XFILL_43_DFFSR_51 gnd vdd FILL
XFILL_63_DFFSR_103 gnd vdd FILL
XFILL_2_MUX2X1_27 gnd vdd FILL
XFILL_63_DFFSR_114 gnd vdd FILL
XFILL_43_DFFSR_62 gnd vdd FILL
XFILL_2_MUX2X1_38 gnd vdd FILL
XFILL_43_DFFSR_73 gnd vdd FILL
XFILL_2_MUX2X1_49 gnd vdd FILL
XFILL_63_DFFSR_125 gnd vdd FILL
XFILL_63_DFFSR_136 gnd vdd FILL
XFILL_43_DFFSR_84 gnd vdd FILL
XFILL_43_DFFSR_95 gnd vdd FILL
XFILL_10_NAND3X1_102 gnd vdd FILL
XFILL_63_DFFSR_147 gnd vdd FILL
XFILL_63_DFFSR_158 gnd vdd FILL
XFILL_10_NAND3X1_113 gnd vdd FILL
XFILL_9_DFFSR_270 gnd vdd FILL
XFILL_10_NAND3X1_124 gnd vdd FILL
XFILL_23_5_2 gnd vdd FILL
XFILL_63_DFFSR_169 gnd vdd FILL
XFILL_6_MUX2X1_15 gnd vdd FILL
XFILL_67_DFFSR_102 gnd vdd FILL
XFILL_22_0_1 gnd vdd FILL
XFILL_6_MUX2X1_26 gnd vdd FILL
XFILL_83_DFFSR_50 gnd vdd FILL
XFILL_6_MUX2X1_37 gnd vdd FILL
XFILL_67_DFFSR_113 gnd vdd FILL
XFILL_83_DFFSR_61 gnd vdd FILL
XFILL_6_MUX2X1_48 gnd vdd FILL
XFILL_8_NOR2X1_109 gnd vdd FILL
XFILL_83_DFFSR_72 gnd vdd FILL
XFILL_83_DFFSR_83 gnd vdd FILL
XFILL_67_DFFSR_124 gnd vdd FILL
XFILL_6_MUX2X1_59 gnd vdd FILL
XFILL_67_DFFSR_135 gnd vdd FILL
XFILL_67_DFFSR_146 gnd vdd FILL
XFILL_10_OAI21X1_3 gnd vdd FILL
XFILL_14_NAND3X1_11 gnd vdd FILL
XFILL_83_DFFSR_94 gnd vdd FILL
XFILL_12_DFFSR_50 gnd vdd FILL
XFILL_67_DFFSR_157 gnd vdd FILL
XFILL_14_NAND3X1_22 gnd vdd FILL
XFILL_12_DFFSR_61 gnd vdd FILL
XFILL_67_DFFSR_168 gnd vdd FILL
XFILL_14_NAND3X1_33 gnd vdd FILL
XFILL_1_MUX2X1_180 gnd vdd FILL
XFILL_12_DFFSR_72 gnd vdd FILL
XFILL_12_DFFSR_83 gnd vdd FILL
XFILL_13_BUFX4_8 gnd vdd FILL
XFILL_1_MUX2X1_191 gnd vdd FILL
XFILL_67_DFFSR_179 gnd vdd FILL
XFILL_14_NAND3X1_44 gnd vdd FILL
XFILL_14_NAND3X1_55 gnd vdd FILL
XFILL_12_DFFSR_94 gnd vdd FILL
XFILL_34_CLKBUF1_11 gnd vdd FILL
XFILL_14_NAND3X1_66 gnd vdd FILL
XFILL_34_CLKBUF1_22 gnd vdd FILL
XFILL_14_NAND3X1_77 gnd vdd FILL
XFILL_23_NOR3X1_2 gnd vdd FILL
XFILL_14_NAND3X1_88 gnd vdd FILL
XFILL_34_CLKBUF1_33 gnd vdd FILL
XFILL_14_OAI21X1_2 gnd vdd FILL
XFILL_14_NAND3X1_99 gnd vdd FILL
XFILL_1_NAND3X1_107 gnd vdd FILL
XFILL_1_NAND3X1_118 gnd vdd FILL
XFILL_52_DFFSR_60 gnd vdd FILL
XFILL_52_DFFSR_71 gnd vdd FILL
XFILL_52_DFFSR_82 gnd vdd FILL
XFILL_11_NOR2X1_60 gnd vdd FILL
XFILL_1_NAND3X1_129 gnd vdd FILL
XFILL_52_DFFSR_93 gnd vdd FILL
XFILL_11_NOR2X1_71 gnd vdd FILL
XFILL_11_NOR2X1_82 gnd vdd FILL
XFILL_2_INVX1_220 gnd vdd FILL
XFILL_11_NOR2X1_93 gnd vdd FILL
XFILL_22_MUX2X1_13 gnd vdd FILL
XFILL_21_DFFSR_70 gnd vdd FILL
XFILL_22_MUX2X1_24 gnd vdd FILL
XFILL_22_MUX2X1_35 gnd vdd FILL
XFILL_21_DFFSR_81 gnd vdd FILL
XFILL_21_DFFSR_92 gnd vdd FILL
XFILL_6_6_2 gnd vdd FILL
XFILL_22_MUX2X1_46 gnd vdd FILL
XFILL_6_NOR3X1_3 gnd vdd FILL
XFILL_22_MUX2X1_57 gnd vdd FILL
XFILL_5_OAI22X1_18 gnd vdd FILL
XFILL_22_MUX2X1_68 gnd vdd FILL
XFILL_5_1_1 gnd vdd FILL
XFILL_5_OAI22X1_29 gnd vdd FILL
XFILL_22_MUX2X1_79 gnd vdd FILL
XFILL_52_DFFSR_190 gnd vdd FILL
XFILL_18_AOI22X1_11 gnd vdd FILL
XFILL_61_DFFSR_80 gnd vdd FILL
XFILL_61_DFFSR_91 gnd vdd FILL
XFILL_4_NAND3X1_50 gnd vdd FILL
XFILL_4_NAND3X1_61 gnd vdd FILL
XFILL_4_NAND3X1_72 gnd vdd FILL
XFILL_8_NAND2X1_30 gnd vdd FILL
XFILL_30_DFFSR_103 gnd vdd FILL
XFILL_8_NAND2X1_41 gnd vdd FILL
XFILL_4_NAND3X1_83 gnd vdd FILL
XFILL_36_DFFSR_2 gnd vdd FILL
XFILL_4_NAND3X1_94 gnd vdd FILL
XFILL_8_NAND2X1_52 gnd vdd FILL
XFILL_30_DFFSR_114 gnd vdd FILL
XFILL_14_5_2 gnd vdd FILL
XFILL_4_DFFSR_60 gnd vdd FILL
XFILL_8_NAND2X1_63 gnd vdd FILL
XFILL_4_DFFSR_71 gnd vdd FILL
XFILL_30_DFFSR_125 gnd vdd FILL
XFILL_30_DFFSR_136 gnd vdd FILL
XFILL_4_DFFSR_82 gnd vdd FILL
XFILL_8_NAND2X1_74 gnd vdd FILL
XFILL_4_DFFSR_93 gnd vdd FILL
XFILL_13_0_1 gnd vdd FILL
XFILL_8_NAND2X1_85 gnd vdd FILL
XFILL_30_DFFSR_147 gnd vdd FILL
XFILL_30_DFFSR_158 gnd vdd FILL
XFILL_8_NAND2X1_96 gnd vdd FILL
XFILL_30_DFFSR_90 gnd vdd FILL
XFILL_30_DFFSR_169 gnd vdd FILL
XFILL_34_DFFSR_102 gnd vdd FILL
XFILL_16_CLKBUF1_16 gnd vdd FILL
XFILL_34_DFFSR_113 gnd vdd FILL
XFILL_11_NAND2X1_4 gnd vdd FILL
XFILL_34_DFFSR_124 gnd vdd FILL
XFILL_16_CLKBUF1_27 gnd vdd FILL
XFILL_16_CLKBUF1_38 gnd vdd FILL
XFILL_34_DFFSR_135 gnd vdd FILL
XFILL_34_DFFSR_146 gnd vdd FILL
XFILL_11_AOI21X1_13 gnd vdd FILL
XFILL_34_DFFSR_157 gnd vdd FILL
XFILL_3_DFFSR_170 gnd vdd FILL
XFILL_34_DFFSR_168 gnd vdd FILL
XFILL_11_AOI21X1_24 gnd vdd FILL
XFILL_11_AOI21X1_35 gnd vdd FILL
XFILL_3_DFFSR_181 gnd vdd FILL
XFILL_11_AOI21X1_46 gnd vdd FILL
XFILL_34_DFFSR_179 gnd vdd FILL
XAND2X2_4 AND2X2_4/A BUFX4_7/Y gnd AND2X2_4/Y vdd AND2X2
XFILL_3_DFFSR_192 gnd vdd FILL
XFILL_38_DFFSR_101 gnd vdd FILL
XFILL_11_AOI21X1_57 gnd vdd FILL
XFILL_11_AOI21X1_68 gnd vdd FILL
XFILL_20_DFFSR_8 gnd vdd FILL
XFILL_38_DFFSR_112 gnd vdd FILL
XFILL_38_DFFSR_123 gnd vdd FILL
XFILL_11_AOI21X1_79 gnd vdd FILL
XFILL_38_DFFSR_134 gnd vdd FILL
XFILL_38_DFFSR_145 gnd vdd FILL
XFILL_38_DFFSR_156 gnd vdd FILL
XFILL_7_DFFSR_180 gnd vdd FILL
XFILL_58_DFFSR_6 gnd vdd FILL
XFILL_38_DFFSR_167 gnd vdd FILL
XFILL_38_DFFSR_178 gnd vdd FILL
XFILL_30_NOR3X1_14 gnd vdd FILL
XFILL_7_DFFSR_191 gnd vdd FILL
XFILL_38_DFFSR_189 gnd vdd FILL
XFILL_30_NOR3X1_25 gnd vdd FILL
XFILL_30_NOR3X1_36 gnd vdd FILL
XFILL_30_NOR3X1_47 gnd vdd FILL
XFILL_80_DFFSR_203 gnd vdd FILL
XFILL_80_DFFSR_214 gnd vdd FILL
XFILL_2_4 gnd vdd FILL
XFILL_80_DFFSR_225 gnd vdd FILL
XFILL_80_DFFSR_236 gnd vdd FILL
XFILL_80_DFFSR_247 gnd vdd FILL
XFILL_80_DFFSR_258 gnd vdd FILL
XFILL_80_DFFSR_269 gnd vdd FILL
XFILL_84_DFFSR_202 gnd vdd FILL
XFILL_84_DFFSR_213 gnd vdd FILL
XFILL_23_CLKBUF1_40 gnd vdd FILL
XFILL_84_DFFSR_224 gnd vdd FILL
XFILL_84_DFFSR_235 gnd vdd FILL
XFILL_11_AOI21X1_9 gnd vdd FILL
XFILL_84_DFFSR_246 gnd vdd FILL
XFILL_64_4_2 gnd vdd FILL
XFILL_6_CLKBUF1_11 gnd vdd FILL
XFILL_84_DFFSR_257 gnd vdd FILL
XFILL_6_CLKBUF1_22 gnd vdd FILL
XFILL_84_DFFSR_268 gnd vdd FILL
XFILL_44_4 gnd vdd FILL
XFILL_6_CLKBUF1_33 gnd vdd FILL
XFILL_0_INVX1_130 gnd vdd FILL
XFILL_14_MUX2X1_107 gnd vdd FILL
XFILL_14_MUX2X1_118 gnd vdd FILL
XFILL_0_INVX1_141 gnd vdd FILL
XFILL_0_INVX1_152 gnd vdd FILL
XFILL_1_AOI21X1_30 gnd vdd FILL
XFILL_14_MUX2X1_129 gnd vdd FILL
XFILL_15_AOI21X1_8 gnd vdd FILL
XFILL_0_INVX1_163 gnd vdd FILL
XFILL_1_AOI21X1_41 gnd vdd FILL
XFILL_1_AOI21X1_52 gnd vdd FILL
XFILL_11_OAI22X1_10 gnd vdd FILL
XFILL_0_INVX1_174 gnd vdd FILL
XFILL_0_INVX1_185 gnd vdd FILL
XFILL_1_AOI21X1_63 gnd vdd FILL
XFILL_11_OAI22X1_21 gnd vdd FILL
XFILL_1_AOI21X1_74 gnd vdd FILL
XFILL_0_INVX1_196 gnd vdd FILL
XFILL_11_OAI22X1_32 gnd vdd FILL
XFILL_11_OAI22X1_43 gnd vdd FILL
XFILL_4_INVX1_140 gnd vdd FILL
XFILL_15_OAI21X1_12 gnd vdd FILL
XFILL_4_INVX1_151 gnd vdd FILL
XFILL_15_OAI21X1_23 gnd vdd FILL
XFILL_4_INVX1_162 gnd vdd FILL
XFILL_15_OAI21X1_34 gnd vdd FILL
XFILL_4_NOR2X1_140 gnd vdd FILL
XFILL_15_OAI21X1_45 gnd vdd FILL
XFILL_4_INVX1_173 gnd vdd FILL
XFILL_4_NOR2X1_151 gnd vdd FILL
XFILL_4_NOR2X1_162 gnd vdd FILL
XFILL_4_INVX1_184 gnd vdd FILL
XFILL_4_NOR2X1_173 gnd vdd FILL
XFILL_4_INVX1_195 gnd vdd FILL
XFILL_4_NOR2X1_184 gnd vdd FILL
XFILL_4_NOR2X1_195 gnd vdd FILL
XFILL_21_MUX2X1_120 gnd vdd FILL
XFILL_2_OAI22X1_2 gnd vdd FILL
XFILL_21_MUX2X1_131 gnd vdd FILL
XFILL_21_MUX2X1_142 gnd vdd FILL
XFILL_21_MUX2X1_153 gnd vdd FILL
XFILL_60_12 gnd vdd FILL
XFILL_21_MUX2X1_164 gnd vdd FILL
XFILL_21_MUX2X1_175 gnd vdd FILL
XFILL_4_MUX2X1_102 gnd vdd FILL
XFILL_4_MUX2X1_113 gnd vdd FILL
XFILL_4_MUX2X1_124 gnd vdd FILL
XFILL_21_MUX2X1_186 gnd vdd FILL
XFILL_4_MUX2X1_135 gnd vdd FILL
XFILL_4_MUX2X1_146 gnd vdd FILL
XFILL_6_OAI22X1_1 gnd vdd FILL
XFILL_4_MUX2X1_157 gnd vdd FILL
XFILL_4_MUX2X1_168 gnd vdd FILL
XFILL_4_MUX2X1_179 gnd vdd FILL
XFILL_51_DFFSR_202 gnd vdd FILL
XFILL_55_4_2 gnd vdd FILL
XFILL_51_DFFSR_213 gnd vdd FILL
XFILL_5_OAI21X1_40 gnd vdd FILL
XFILL_51_DFFSR_224 gnd vdd FILL
XFILL_51_DFFSR_235 gnd vdd FILL
XFILL_51_DFFSR_246 gnd vdd FILL
XFILL_75_DFFSR_19 gnd vdd FILL
XFILL_51_DFFSR_257 gnd vdd FILL
XFILL_51_DFFSR_268 gnd vdd FILL
XFILL_5_DFFSR_1 gnd vdd FILL
XFILL_55_DFFSR_201 gnd vdd FILL
XFILL_18_MUX2X1_9 gnd vdd FILL
XFILL_55_DFFSR_212 gnd vdd FILL
XFILL_55_DFFSR_223 gnd vdd FILL
XFILL_55_DFFSR_234 gnd vdd FILL
XFILL_11_NAND3X1_103 gnd vdd FILL
XFILL_9_BUFX4_20 gnd vdd FILL
XFILL_11_NAND3X1_114 gnd vdd FILL
XFILL_55_DFFSR_245 gnd vdd FILL
XFILL_11_NAND3X1_125 gnd vdd FILL
XFILL_55_DFFSR_256 gnd vdd FILL
XFILL_9_BUFX4_31 gnd vdd FILL
XFILL_55_DFFSR_267 gnd vdd FILL
XFILL_9_BUFX4_42 gnd vdd FILL
XFILL_10_CLKBUF1_8 gnd vdd FILL
XFILL_82_DFFSR_101 gnd vdd FILL
XFILL_9_BUFX4_53 gnd vdd FILL
XFILL_9_BUFX4_64 gnd vdd FILL
XFILL_59_DFFSR_200 gnd vdd FILL
XFILL_82_DFFSR_112 gnd vdd FILL
XFILL_59_DFFSR_211 gnd vdd FILL
XFILL_44_DFFSR_18 gnd vdd FILL
XFILL_9_BUFX4_75 gnd vdd FILL
XFILL_0_BUFX2_7 gnd vdd FILL
XFILL_59_DFFSR_222 gnd vdd FILL
XFILL_44_DFFSR_29 gnd vdd FILL
XFILL_82_DFFSR_123 gnd vdd FILL
XFILL_82_DFFSR_134 gnd vdd FILL
XFILL_59_DFFSR_233 gnd vdd FILL
XFILL_9_BUFX4_86 gnd vdd FILL
XFILL_9_BUFX4_97 gnd vdd FILL
XFILL_82_DFFSR_145 gnd vdd FILL
XFILL_59_DFFSR_244 gnd vdd FILL
XFILL_82_DFFSR_156 gnd vdd FILL
XFILL_59_DFFSR_255 gnd vdd FILL
XFILL_82_DFFSR_167 gnd vdd FILL
XFILL_59_DFFSR_266 gnd vdd FILL
XFILL_14_CLKBUF1_7 gnd vdd FILL
XFILL_82_DFFSR_178 gnd vdd FILL
XFILL_86_DFFSR_100 gnd vdd FILL
XFILL_82_DFFSR_189 gnd vdd FILL
XFILL_2_DFFSR_204 gnd vdd FILL
XFILL_2_DFFSR_215 gnd vdd FILL
XFILL_84_DFFSR_17 gnd vdd FILL
XFILL_86_DFFSR_111 gnd vdd FILL
XFILL_2_DFFSR_226 gnd vdd FILL
XFILL_86_DFFSR_122 gnd vdd FILL
XFILL_7_NAND3X1_16 gnd vdd FILL
XFILL_84_DFFSR_28 gnd vdd FILL
XFILL_86_DFFSR_133 gnd vdd FILL
XFILL_2_DFFSR_237 gnd vdd FILL
XFILL_84_DFFSR_39 gnd vdd FILL
XFILL_7_NAND3X1_27 gnd vdd FILL
XFILL_86_DFFSR_144 gnd vdd FILL
XFILL_2_NAND3X1_108 gnd vdd FILL
XFILL_2_DFFSR_248 gnd vdd FILL
XFILL_7_NAND3X1_38 gnd vdd FILL
XFILL_86_DFFSR_155 gnd vdd FILL
XFILL_10_BUFX4_102 gnd vdd FILL
XFILL_13_DFFSR_17 gnd vdd FILL
XFILL_2_NAND3X1_119 gnd vdd FILL
XFILL_7_NAND3X1_49 gnd vdd FILL
XFILL_2_DFFSR_259 gnd vdd FILL
XFILL_86_DFFSR_166 gnd vdd FILL
XFILL_86_DFFSR_177 gnd vdd FILL
XFILL_13_DFFSR_28 gnd vdd FILL
XFILL_13_DFFSR_39 gnd vdd FILL
XFILL_18_CLKBUF1_6 gnd vdd FILL
XFILL_3_NAND3X1_3 gnd vdd FILL
XFILL_86_DFFSR_188 gnd vdd FILL
XFILL_6_DFFSR_203 gnd vdd FILL
XFILL_86_DFFSR_199 gnd vdd FILL
XFILL_6_DFFSR_214 gnd vdd FILL
XFILL_11_OR2X2_1 gnd vdd FILL
XFILL_6_DFFSR_225 gnd vdd FILL
XFILL_6_DFFSR_236 gnd vdd FILL
XFILL_6_DFFSR_247 gnd vdd FILL
XFILL_14_BUFX4_101 gnd vdd FILL
XFILL_53_DFFSR_16 gnd vdd FILL
XFILL_6_DFFSR_258 gnd vdd FILL
XFILL_6_DFFSR_269 gnd vdd FILL
XFILL_53_DFFSR_27 gnd vdd FILL
XFILL_53_DFFSR_38 gnd vdd FILL
XFILL_53_DFFSR_49 gnd vdd FILL
XFILL_7_NAND3X1_2 gnd vdd FILL
XMUX2X1_16 MUX2X1_66/A INVX1_29/Y MUX2X1_16/S gnd DFFSR_27/D vdd MUX2X1
XFILL_0_NAND2X1_18 gnd vdd FILL
XFILL_46_4_2 gnd vdd FILL
XMUX2X1_27 BUFX4_71/Y INVX1_40/Y NOR2X1_12/B gnd MUX2X1_27/Y vdd MUX2X1
XFILL_0_NAND2X1_29 gnd vdd FILL
XMUX2X1_38 INVX1_51/Y BUFX4_66/Y NAND2X1_5/Y gnd MUX2X1_38/Y vdd MUX2X1
XFILL_24_DFFSR_9 gnd vdd FILL
XMUX2X1_49 INVX1_62/Y MUX2X1_7/B NAND2X1_7/Y gnd MUX2X1_49/Y vdd MUX2X1
XFILL_22_DFFSR_15 gnd vdd FILL
XFILL_22_DFFSR_26 gnd vdd FILL
XFILL_22_DFFSR_37 gnd vdd FILL
XFILL_13_BUFX4_80 gnd vdd FILL
XFILL_22_DFFSR_48 gnd vdd FILL
XFILL_22_DFFSR_59 gnd vdd FILL
XFILL_13_BUFX4_91 gnd vdd FILL
XFILL_10_MUX2X1_160 gnd vdd FILL
XFILL_10_MUX2X1_171 gnd vdd FILL
XFILL_23_9 gnd vdd FILL
XFILL_62_DFFSR_14 gnd vdd FILL
XFILL_10_MUX2X1_182 gnd vdd FILL
XFILL_22_DFFSR_201 gnd vdd FILL
XFILL_62_DFFSR_25 gnd vdd FILL
XFILL_10_MUX2X1_193 gnd vdd FILL
XFILL_62_DFFSR_36 gnd vdd FILL
XFILL_22_DFFSR_212 gnd vdd FILL
XFILL_22_DFFSR_223 gnd vdd FILL
XFILL_62_DFFSR_47 gnd vdd FILL
XFILL_22_DFFSR_234 gnd vdd FILL
XFILL_16_8 gnd vdd FILL
XFILL_3_AOI22X1_8 gnd vdd FILL
XFILL_62_DFFSR_58 gnd vdd FILL
XFILL_62_DFFSR_69 gnd vdd FILL
XFILL_22_DFFSR_245 gnd vdd FILL
XFILL_22_DFFSR_256 gnd vdd FILL
XFILL_22_DFFSR_267 gnd vdd FILL
XFILL_3_INVX1_207 gnd vdd FILL
XFILL_26_DFFSR_200 gnd vdd FILL
XFILL_3_INVX1_218 gnd vdd FILL
XFILL_26_CLKBUF1_17 gnd vdd FILL
XFILL_26_CLKBUF1_28 gnd vdd FILL
XFILL_26_DFFSR_211 gnd vdd FILL
XFILL_5_DFFSR_16 gnd vdd FILL
XFILL_26_DFFSR_222 gnd vdd FILL
XDFFSR_8 DFFSR_8/Q DFFSR_8/CLK DFFSR_8/R vdd DFFSR_8/D gnd vdd DFFSR
XFILL_5_DFFSR_27 gnd vdd FILL
XFILL_26_DFFSR_233 gnd vdd FILL
XFILL_5_DFFSR_38 gnd vdd FILL
XFILL_7_AOI22X1_7 gnd vdd FILL
XFILL_26_CLKBUF1_39 gnd vdd FILL
XFILL_31_DFFSR_13 gnd vdd FILL
XFILL_26_DFFSR_244 gnd vdd FILL
XFILL_31_DFFSR_24 gnd vdd FILL
XFILL_5_DFFSR_49 gnd vdd FILL
XFILL_31_DFFSR_35 gnd vdd FILL
XFILL_26_DFFSR_255 gnd vdd FILL
XFILL_31_DFFSR_46 gnd vdd FILL
XFILL_26_DFFSR_266 gnd vdd FILL
XFILL_31_DFFSR_57 gnd vdd FILL
XFILL_7_INVX1_206 gnd vdd FILL
XINVX1_220 DFFSR_63/Q gnd INVX1_220/Y vdd INVX1
XFILL_53_DFFSR_100 gnd vdd FILL
XFILL_31_DFFSR_68 gnd vdd FILL
XFILL_53_DFFSR_111 gnd vdd FILL
XFILL_7_INVX1_217 gnd vdd FILL
XFILL_31_DFFSR_79 gnd vdd FILL
XFILL_7_INVX1_70 gnd vdd FILL
XFILL_7_INVX1_228 gnd vdd FILL
XFILL_53_DFFSR_122 gnd vdd FILL
XFILL_4_AOI21X1_18 gnd vdd FILL
XFILL_7_INVX1_81 gnd vdd FILL
XFILL_7_INVX1_92 gnd vdd FILL
XFILL_53_DFFSR_133 gnd vdd FILL
XFILL_71_DFFSR_12 gnd vdd FILL
XFILL_4_AOI21X1_29 gnd vdd FILL
XFILL_53_DFFSR_144 gnd vdd FILL
XFILL_53_DFFSR_155 gnd vdd FILL
XFILL_71_DFFSR_23 gnd vdd FILL
XFILL_71_DFFSR_34 gnd vdd FILL
XFILL_53_DFFSR_166 gnd vdd FILL
XFILL_14_MUX2X1_2 gnd vdd FILL
XFILL_71_DFFSR_45 gnd vdd FILL
XFILL_71_DFFSR_56 gnd vdd FILL
XFILL_53_DFFSR_177 gnd vdd FILL
XFILL_71_DFFSR_67 gnd vdd FILL
XFILL_53_DFFSR_188 gnd vdd FILL
XFILL_57_DFFSR_110 gnd vdd FILL
XFILL_53_DFFSR_199 gnd vdd FILL
XFILL_7_NOR2X1_106 gnd vdd FILL
XFILL_71_DFFSR_78 gnd vdd FILL
XFILL_57_DFFSR_121 gnd vdd FILL
XFILL_71_DFFSR_89 gnd vdd FILL
XFILL_7_NOR2X1_117 gnd vdd FILL
XFILL_57_DFFSR_132 gnd vdd FILL
XFILL_7_NOR2X1_128 gnd vdd FILL
XFILL_57_DFFSR_143 gnd vdd FILL
XFILL_57_DFFSR_154 gnd vdd FILL
XFILL_7_NOR2X1_139 gnd vdd FILL
XNAND2X1_20 BUFX4_58/Y NOR2X1_30/Y gnd OAI22X1_33/B vdd NAND2X1
XFILL_57_DFFSR_165 gnd vdd FILL
XFILL_13_NAND3X1_30 gnd vdd FILL
XNAND2X1_31 BUFX4_1/Y AND2X2_4/A gnd OAI22X1_48/D vdd NAND2X1
XFILL_13_NAND3X1_41 gnd vdd FILL
XFILL_57_DFFSR_176 gnd vdd FILL
XFILL_40_DFFSR_11 gnd vdd FILL
XNAND2X1_42 BUFX4_6/Y NOR3X1_51/Y gnd NOR2X1_80/B vdd NAND2X1
XFILL_0_DFFSR_103 gnd vdd FILL
XNAND2X1_53 BUFX4_92/Y NOR2X1_31/Y gnd OAI22X1_4/B vdd NAND2X1
XFILL_57_DFFSR_187 gnd vdd FILL
XFILL_40_DFFSR_22 gnd vdd FILL
XFILL_0_DFFSR_114 gnd vdd FILL
XFILL_13_NAND3X1_52 gnd vdd FILL
XFILL_57_DFFSR_198 gnd vdd FILL
XNAND2X1_64 INVX2_2/A NOR2X1_38/Y gnd NOR2X1_86/B vdd NAND2X1
XFILL_13_NAND3X1_63 gnd vdd FILL
XFILL_65_7_0 gnd vdd FILL
XFILL_13_NAND3X1_74 gnd vdd FILL
XFILL_5_BUFX4_90 gnd vdd FILL
XNAND2X1_75 NOR2X1_100/Y NOR2X1_99/Y gnd NOR3X1_43/B vdd NAND2X1
XFILL_40_DFFSR_33 gnd vdd FILL
XFILL_0_DFFSR_125 gnd vdd FILL
XFILL_0_DFFSR_136 gnd vdd FILL
XFILL_33_CLKBUF1_30 gnd vdd FILL
XFILL_11_NOR3X1_8 gnd vdd FILL
XFILL_13_NAND3X1_85 gnd vdd FILL
XNAND2X1_86 AOI22X1_1/A AOI22X1_1/B gnd AND2X2_2/A vdd NAND2X1
XFILL_40_DFFSR_44 gnd vdd FILL
XFILL_40_DFFSR_55 gnd vdd FILL
XFILL_13_NAND3X1_96 gnd vdd FILL
XFILL_37_4_2 gnd vdd FILL
XFILL_0_DFFSR_147 gnd vdd FILL
XFILL_33_CLKBUF1_41 gnd vdd FILL
XFILL_0_DFFSR_158 gnd vdd FILL
XFILL_40_DFFSR_66 gnd vdd FILL
XFILL_40_DFFSR_77 gnd vdd FILL
XFILL_42_1 gnd vdd FILL
XFILL_0_DFFSR_169 gnd vdd FILL
XFILL_40_DFFSR_88 gnd vdd FILL
XFILL_4_DFFSR_102 gnd vdd FILL
XFILL_40_DFFSR_99 gnd vdd FILL
XFILL_80_DFFSR_10 gnd vdd FILL
XFILL_80_DFFSR_21 gnd vdd FILL
XFILL_4_DFFSR_113 gnd vdd FILL
XFILL_80_DFFSR_32 gnd vdd FILL
XFILL_4_DFFSR_124 gnd vdd FILL
XFILL_80_DFFSR_43 gnd vdd FILL
XFILL_4_DFFSR_135 gnd vdd FILL
XFILL_4_DFFSR_146 gnd vdd FILL
XFILL_80_DFFSR_54 gnd vdd FILL
XFILL_4_DFFSR_157 gnd vdd FILL
XFILL_80_DFFSR_65 gnd vdd FILL
XFILL_80_DFFSR_76 gnd vdd FILL
XFILL_4_DFFSR_168 gnd vdd FILL
XFILL_80_DFFSR_87 gnd vdd FILL
XFILL_4_DFFSR_179 gnd vdd FILL
XFILL_80_DFFSR_98 gnd vdd FILL
XFILL_8_DFFSR_101 gnd vdd FILL
XFILL_7_NOR2X1_3 gnd vdd FILL
XFILL_12_MUX2X1_10 gnd vdd FILL
XFILL_8_DFFSR_112 gnd vdd FILL
XFILL_12_MUX2X1_21 gnd vdd FILL
XFILL_8_DFFSR_123 gnd vdd FILL
XFILL_8_DFFSR_134 gnd vdd FILL
XFILL_12_MUX2X1_32 gnd vdd FILL
XFILL_8_DFFSR_145 gnd vdd FILL
XFILL_20_3_2 gnd vdd FILL
XFILL_12_MUX2X1_43 gnd vdd FILL
XFILL_8_DFFSR_156 gnd vdd FILL
XFILL_12_MUX2X1_54 gnd vdd FILL
XFILL_4_OAI22X1_15 gnd vdd FILL
XFILL_8_DFFSR_167 gnd vdd FILL
XFILL_12_MUX2X1_65 gnd vdd FILL
XFILL_8_DFFSR_178 gnd vdd FILL
XFILL_12_MUX2X1_76 gnd vdd FILL
XFILL_20_NOR3X1_6 gnd vdd FILL
XFILL_4_OAI22X1_26 gnd vdd FILL
XFILL_0_NOR3X1_14 gnd vdd FILL
XFILL_4_OAI22X1_37 gnd vdd FILL
XFILL_12_MUX2X1_87 gnd vdd FILL
XFILL_8_DFFSR_189 gnd vdd FILL
XFILL_0_NOR3X1_25 gnd vdd FILL
XFILL_0_NOR3X1_36 gnd vdd FILL
XFILL_12_MUX2X1_98 gnd vdd FILL
XFILL_4_OAI22X1_48 gnd vdd FILL
XFILL_8_OAI21X1_17 gnd vdd FILL
XFILL_16_MUX2X1_20 gnd vdd FILL
XFILL_0_NOR3X1_47 gnd vdd FILL
XFILL_16_MUX2X1_31 gnd vdd FILL
XFILL_8_OAI21X1_28 gnd vdd FILL
XFILL_16_MUX2X1_42 gnd vdd FILL
XFILL_8_OAI21X1_39 gnd vdd FILL
XFILL_16_MUX2X1_53 gnd vdd FILL
XFILL_6_MUX2X1_1 gnd vdd FILL
XFILL_16_MUX2X1_64 gnd vdd FILL
XFILL_16_MUX2X1_75 gnd vdd FILL
XFILL_4_NOR3X1_13 gnd vdd FILL
XFILL_16_MUX2X1_86 gnd vdd FILL
XFILL_4_NOR3X1_24 gnd vdd FILL
XFILL_41_DFFSR_3 gnd vdd FILL
XFILL_16_MUX2X1_97 gnd vdd FILL
XFILL_4_NOR3X1_35 gnd vdd FILL
XFILL_4_NOR3X1_46 gnd vdd FILL
XFILL_20_DFFSR_100 gnd vdd FILL
XFILL_3_NAND3X1_80 gnd vdd FILL
XFILL_9_DFFSR_2 gnd vdd FILL
XFILL_3_NAND3X1_91 gnd vdd FILL
XFILL_20_DFFSR_111 gnd vdd FILL
XFILL_7_NAND2X1_60 gnd vdd FILL
XFILL_1_NOR2X1_206 gnd vdd FILL
XFILL_20_DFFSR_122 gnd vdd FILL
XFILL_20_DFFSR_133 gnd vdd FILL
XFILL_79_DFFSR_1 gnd vdd FILL
XFILL_7_NAND2X1_71 gnd vdd FILL
XFILL_20_DFFSR_144 gnd vdd FILL
XFILL_7_NAND2X1_82 gnd vdd FILL
XFILL_20_DFFSR_155 gnd vdd FILL
XFILL_7_NAND2X1_93 gnd vdd FILL
XFILL_8_NOR3X1_12 gnd vdd FILL
XFILL_20_DFFSR_166 gnd vdd FILL
XFILL_8_NOR3X1_23 gnd vdd FILL
XFILL_3_NOR3X1_7 gnd vdd FILL
XFILL_8_NOR3X1_34 gnd vdd FILL
XFILL_20_DFFSR_177 gnd vdd FILL
XFILL_1_INVX1_106 gnd vdd FILL
XFILL_1_INVX1_117 gnd vdd FILL
XFILL_20_DFFSR_188 gnd vdd FILL
XFILL_8_NOR3X1_45 gnd vdd FILL
XFILL_24_DFFSR_110 gnd vdd FILL
XFILL_20_DFFSR_199 gnd vdd FILL
XFILL_15_CLKBUF1_13 gnd vdd FILL
XFILL_15_CLKBUF1_24 gnd vdd FILL
XFILL_1_INVX1_128 gnd vdd FILL
XFILL_24_DFFSR_121 gnd vdd FILL
XFILL_4_BUFX2_8 gnd vdd FILL
XFILL_1_INVX1_139 gnd vdd FILL
XFILL_24_DFFSR_132 gnd vdd FILL
XFILL_15_CLKBUF1_35 gnd vdd FILL
XFILL_24_DFFSR_143 gnd vdd FILL
XFILL_10_AOI21X1_10 gnd vdd FILL
XFILL_24_DFFSR_154 gnd vdd FILL
XFILL_10_AOI21X1_21 gnd vdd FILL
XFILL_24_DFFSR_165 gnd vdd FILL
XFILL_56_7_0 gnd vdd FILL
XFILL_10_AOI21X1_32 gnd vdd FILL
XFILL_24_DFFSR_176 gnd vdd FILL
XFILL_10_AOI21X1_43 gnd vdd FILL
XFILL_5_INVX1_105 gnd vdd FILL
XFILL_28_4_2 gnd vdd FILL
XFILL_5_INVX1_116 gnd vdd FILL
XFILL_24_DFFSR_187 gnd vdd FILL
XFILL_10_AOI21X1_54 gnd vdd FILL
XFILL_3_4_2 gnd vdd FILL
XFILL_24_DFFSR_198 gnd vdd FILL
XFILL_1_DFFSR_20 gnd vdd FILL
XFILL_10_AOI21X1_65 gnd vdd FILL
XFILL_5_INVX1_127 gnd vdd FILL
XFILL_28_DFFSR_120 gnd vdd FILL
XFILL_1_DFFSR_31 gnd vdd FILL
XFILL_10_AOI21X1_76 gnd vdd FILL
XFILL_28_DFFSR_131 gnd vdd FILL
XFILL_1_DFFSR_42 gnd vdd FILL
XFILL_5_INVX1_138 gnd vdd FILL
XFILL_1_DFFSR_53 gnd vdd FILL
XFILL_5_INVX1_149 gnd vdd FILL
XFILL_28_DFFSR_142 gnd vdd FILL
XFILL_28_DFFSR_153 gnd vdd FILL
XFILL_1_DFFSR_64 gnd vdd FILL
XFILL_63_DFFSR_7 gnd vdd FILL
XFILL_1_DFFSR_75 gnd vdd FILL
XFILL_28_DFFSR_164 gnd vdd FILL
XFILL_28_DFFSR_175 gnd vdd FILL
XFILL_1_DFFSR_86 gnd vdd FILL
XFILL_20_NOR3X1_11 gnd vdd FILL
XFILL_1_DFFSR_97 gnd vdd FILL
XFILL_28_DFFSR_186 gnd vdd FILL
XFILL_20_NOR3X1_22 gnd vdd FILL
XFILL_28_DFFSR_197 gnd vdd FILL
XFILL_20_NOR3X1_33 gnd vdd FILL
XFILL_20_NOR3X1_44 gnd vdd FILL
XFILL_70_DFFSR_200 gnd vdd FILL
XFILL_70_DFFSR_211 gnd vdd FILL
XFILL_70_DFFSR_222 gnd vdd FILL
XFILL_70_DFFSR_233 gnd vdd FILL
XFILL_12_NAND3X1_104 gnd vdd FILL
XFILL_12_NAND3X1_115 gnd vdd FILL
XFILL_70_DFFSR_244 gnd vdd FILL
XFILL_24_NOR3X1_10 gnd vdd FILL
XFILL_70_DFFSR_255 gnd vdd FILL
XFILL_11_3_2 gnd vdd FILL
XFILL_12_NAND3X1_126 gnd vdd FILL
XFILL_70_DFFSR_266 gnd vdd FILL
XFILL_24_NOR3X1_21 gnd vdd FILL
XFILL_24_NOR3X1_32 gnd vdd FILL
XFILL_24_NOR3X1_43 gnd vdd FILL
XFILL_74_DFFSR_210 gnd vdd FILL
XFILL_74_DFFSR_221 gnd vdd FILL
XFILL_74_DFFSR_232 gnd vdd FILL
XFILL_74_DFFSR_243 gnd vdd FILL
XFILL_74_DFFSR_254 gnd vdd FILL
XFILL_3_BUFX4_2 gnd vdd FILL
XFILL_74_DFFSR_265 gnd vdd FILL
XFILL_28_NOR3X1_20 gnd vdd FILL
XFILL_5_CLKBUF1_30 gnd vdd FILL
XFILL_28_NOR3X1_31 gnd vdd FILL
XFILL_5_CLKBUF1_41 gnd vdd FILL
XFILL_28_NOR3X1_42 gnd vdd FILL
XOAI22X1_2 INVX1_89/Y OAI22X1_6/B INVX1_93/Y OAI22X1_6/D gnd OAI22X1_2/Y vdd OAI22X1
XFILL_13_MUX2X1_104 gnd vdd FILL
XFILL_13_MUX2X1_115 gnd vdd FILL
XFILL_13_MUX2X1_126 gnd vdd FILL
XFILL_78_DFFSR_220 gnd vdd FILL
XFILL_78_DFFSR_231 gnd vdd FILL
XFILL_78_DFFSR_242 gnd vdd FILL
XFILL_13_MUX2X1_137 gnd vdd FILL
XFILL_3_NAND3X1_109 gnd vdd FILL
XFILL_13_MUX2X1_148 gnd vdd FILL
XFILL_78_DFFSR_253 gnd vdd FILL
XFILL_13_MUX2X1_159 gnd vdd FILL
XFILL_0_AOI21X1_60 gnd vdd FILL
XFILL_0_AOI21X1_71 gnd vdd FILL
XFILL_78_DFFSR_264 gnd vdd FILL
XFILL_78_DFFSR_275 gnd vdd FILL
XFILL_33_CLKBUF1_5 gnd vdd FILL
XFILL_10_OAI22X1_40 gnd vdd FILL
XFILL_10_OAI22X1_51 gnd vdd FILL
XFILL_14_OAI21X1_20 gnd vdd FILL
XFILL_14_OAI21X1_31 gnd vdd FILL
XFILL_14_OAI21X1_42 gnd vdd FILL
XFILL_3_NOR2X1_170 gnd vdd FILL
XFILL_2_INVX1_6 gnd vdd FILL
XFILL_3_NOR2X1_181 gnd vdd FILL
XFILL_3_NOR2X1_192 gnd vdd FILL
XFILL_47_7_0 gnd vdd FILL
XFILL_19_4_2 gnd vdd FILL
XFILL_61_2_2 gnd vdd FILL
XFILL_20_MUX2X1_150 gnd vdd FILL
XFILL_21_6 gnd vdd FILL
XFILL_20_MUX2X1_161 gnd vdd FILL
XFILL_20_MUX2X1_172 gnd vdd FILL
XFILL_3_MUX2X1_110 gnd vdd FILL
XFILL_20_MUX2X1_183 gnd vdd FILL
XFILL_3_MUX2X1_121 gnd vdd FILL
XFILL_87_DFFSR_109 gnd vdd FILL
XFILL_14_5 gnd vdd FILL
XFILL_20_MUX2X1_194 gnd vdd FILL
XFILL_3_MUX2X1_132 gnd vdd FILL
XFILL_30_6_0 gnd vdd FILL
XFILL_3_MUX2X1_143 gnd vdd FILL
XFILL_14_BUFX4_14 gnd vdd FILL
XFILL_3_MUX2X1_154 gnd vdd FILL
XFILL_14_BUFX4_25 gnd vdd FILL
XFILL_3_MUX2X1_165 gnd vdd FILL
XFILL_14_BUFX4_36 gnd vdd FILL
XFILL_14_BUFX4_47 gnd vdd FILL
XFILL_3_MUX2X1_176 gnd vdd FILL
XFILL_3_MUX2X1_187 gnd vdd FILL
XDFFSR_204 INVX1_95/A CLKBUF1_7/Y BUFX4_21/Y vdd MUX2X1_82/Y gnd vdd DFFSR
XFILL_14_BUFX4_58 gnd vdd FILL
XDFFSR_215 INVX1_82/A CLKBUF1_4/Y DFFSR_57/R vdd MUX2X1_69/Y gnd vdd DFFSR
XFILL_14_BUFX4_69 gnd vdd FILL
XDFFSR_226 INVX1_75/A CLKBUF1_26/Y DFFSR_4/R vdd MUX2X1_62/Y gnd vdd DFFSR
XDFFSR_237 INVX1_60/A CLKBUF1_5/Y BUFX4_23/Y vdd MUX2X1_47/Y gnd vdd DFFSR
XFILL_41_DFFSR_210 gnd vdd FILL
XDFFSR_248 INVX1_53/A DFFSR_39/CLK DFFSR_45/R vdd MUX2X1_40/Y gnd vdd DFFSR
XFILL_41_DFFSR_221 gnd vdd FILL
XDFFSR_259 INVX1_41/A DFFSR_1/CLK BUFX4_54/Y vdd MUX2X1_28/Y gnd vdd DFFSR
XFILL_41_DFFSR_232 gnd vdd FILL
XFILL_41_DFFSR_243 gnd vdd FILL
XFILL_41_DFFSR_254 gnd vdd FILL
XFILL_0_NOR2X1_80 gnd vdd FILL
XFILL_41_DFFSR_265 gnd vdd FILL
XFILL_0_NOR2X1_91 gnd vdd FILL
XFILL_45_DFFSR_220 gnd vdd FILL
XFILL_80_DFFSR_1 gnd vdd FILL
XFILL_45_DFFSR_231 gnd vdd FILL
XFILL_45_DFFSR_242 gnd vdd FILL
XFILL_45_DFFSR_253 gnd vdd FILL
XFILL_45_DFFSR_264 gnd vdd FILL
XFILL_45_DFFSR_275 gnd vdd FILL
XFILL_4_NOR2X1_90 gnd vdd FILL
XFILL_72_DFFSR_120 gnd vdd FILL
XFILL_72_DFFSR_131 gnd vdd FILL
XFILL_49_DFFSR_230 gnd vdd FILL
XFILL_72_DFFSR_142 gnd vdd FILL
XFILL_49_DFFSR_241 gnd vdd FILL
XFILL_9_AND2X2_7 gnd vdd FILL
XFILL_72_DFFSR_153 gnd vdd FILL
XFILL_49_DFFSR_252 gnd vdd FILL
XFILL_38_7_0 gnd vdd FILL
XFILL_72_DFFSR_164 gnd vdd FILL
XFILL_72_DFFSR_175 gnd vdd FILL
XFILL_49_DFFSR_263 gnd vdd FILL
XFILL_49_DFFSR_274 gnd vdd FILL
XFILL_72_DFFSR_186 gnd vdd FILL
XFILL_72_DFFSR_197 gnd vdd FILL
XFILL_6_NAND3X1_13 gnd vdd FILL
XFILL_76_DFFSR_130 gnd vdd FILL
XFILL_6_NAND3X1_24 gnd vdd FILL
XFILL_6_NAND3X1_35 gnd vdd FILL
XFILL_76_DFFSR_141 gnd vdd FILL
XFILL_76_DFFSR_152 gnd vdd FILL
XFILL_6_NAND3X1_46 gnd vdd FILL
XFILL_6_NAND3X1_57 gnd vdd FILL
XFILL_76_DFFSR_163 gnd vdd FILL
XFILL_45_DFFSR_4 gnd vdd FILL
XFILL_76_DFFSR_174 gnd vdd FILL
XFILL_6_NAND3X1_68 gnd vdd FILL
XFILL_6_BUFX4_13 gnd vdd FILL
XFILL_52_2_2 gnd vdd FILL
XFILL_76_DFFSR_185 gnd vdd FILL
XFILL_6_NAND3X1_79 gnd vdd FILL
XFILL_6_BUFX4_24 gnd vdd FILL
XFILL_76_DFFSR_196 gnd vdd FILL
XFILL_6_BUFX4_35 gnd vdd FILL
XFILL_27_DFFSR_209 gnd vdd FILL
XFILL_6_BUFX4_46 gnd vdd FILL
XFILL_6_BUFX4_57 gnd vdd FILL
XFILL_6_BUFX4_68 gnd vdd FILL
XFILL_6_BUFX4_79 gnd vdd FILL
XFILL_21_6_0 gnd vdd FILL
XFILL_0_NAND2X1_2 gnd vdd FILL
XFILL_54_DFFSR_109 gnd vdd FILL
XFILL_8_BUFX2_9 gnd vdd FILL
XFILL_4_NAND2X1_1 gnd vdd FILL
XFILL_58_DFFSR_108 gnd vdd FILL
XFILL_58_DFFSR_119 gnd vdd FILL
XFILL_67_DFFSR_8 gnd vdd FILL
XFILL_13_AND2X2_1 gnd vdd FILL
XFILL_12_DFFSR_220 gnd vdd FILL
XFILL_12_DFFSR_231 gnd vdd FILL
XFILL_12_DFFSR_242 gnd vdd FILL
XFILL_12_DFFSR_253 gnd vdd FILL
XFILL_12_DFFSR_264 gnd vdd FILL
XFILL_12_DFFSR_275 gnd vdd FILL
XFILL_25_CLKBUF1_14 gnd vdd FILL
XFILL_25_CLKBUF1_25 gnd vdd FILL
XFILL_25_CLKBUF1_36 gnd vdd FILL
XFILL_4_7_0 gnd vdd FILL
XFILL_29_7_0 gnd vdd FILL
XFILL_0_AOI21X1_7 gnd vdd FILL
XFILL_10_BUFX4_40 gnd vdd FILL
XFILL_16_DFFSR_230 gnd vdd FILL
XFILL_10_BUFX4_51 gnd vdd FILL
XFILL_16_DFFSR_241 gnd vdd FILL
XFILL_10_BUFX4_62 gnd vdd FILL
XFILL_7_BUFX4_3 gnd vdd FILL
XFILL_10_BUFX4_73 gnd vdd FILL
XFILL_16_DFFSR_252 gnd vdd FILL
XFILL_16_DFFSR_263 gnd vdd FILL
XFILL_16_DFFSR_274 gnd vdd FILL
XFILL_10_BUFX4_84 gnd vdd FILL
XFILL_8_CLKBUF1_18 gnd vdd FILL
XFILL_10_BUFX4_95 gnd vdd FILL
XFILL_8_CLKBUF1_29 gnd vdd FILL
XFILL_13_MUX2X1_19 gnd vdd FILL
XFILL_3_AOI21X1_15 gnd vdd FILL
XFILL_43_DFFSR_130 gnd vdd FILL
XFILL_43_2_2 gnd vdd FILL
XFILL_4_AOI21X1_6 gnd vdd FILL
XFILL_3_AOI21X1_26 gnd vdd FILL
XFILL_3_AOI21X1_37 gnd vdd FILL
XFILL_43_DFFSR_141 gnd vdd FILL
XFILL_43_DFFSR_152 gnd vdd FILL
XFILL_43_DFFSR_163 gnd vdd FILL
XFILL_3_AOI21X1_48 gnd vdd FILL
XFILL_3_AOI21X1_59 gnd vdd FILL
XFILL_43_DFFSR_174 gnd vdd FILL
XFILL_13_OAI22X1_17 gnd vdd FILL
XOAI21X1_18 INVX1_36/Y OAI21X1_9/B OAI21X1_18/C gnd NOR2X1_81/B vdd OAI21X1
XFILL_13_OAI22X1_28 gnd vdd FILL
XOAI21X1_29 INVX1_149/Y OAI21X1_4/B OAI21X1_29/C gnd OAI21X1_29/Y vdd OAI21X1
XFILL_17_MUX2X1_18 gnd vdd FILL
XFILL_43_DFFSR_185 gnd vdd FILL
XFILL_17_MUX2X1_29 gnd vdd FILL
XFILL_13_OAI22X1_39 gnd vdd FILL
XFILL_43_DFFSR_196 gnd vdd FILL
XFILL_6_NOR2X1_103 gnd vdd FILL
XFILL_6_NOR2X1_114 gnd vdd FILL
XFILL_12_6_0 gnd vdd FILL
XFILL_6_NOR2X1_125 gnd vdd FILL
XFILL_8_AOI21X1_5 gnd vdd FILL
XFILL_47_DFFSR_140 gnd vdd FILL
XFILL_6_NOR2X1_136 gnd vdd FILL
XFILL_47_DFFSR_151 gnd vdd FILL
XFILL_47_DFFSR_162 gnd vdd FILL
XFILL_6_NOR2X1_147 gnd vdd FILL
XFILL_13_NAND3X1_105 gnd vdd FILL
XFILL_6_NOR2X1_158 gnd vdd FILL
XFILL_13_NAND3X1_116 gnd vdd FILL
XFILL_47_DFFSR_173 gnd vdd FILL
XFILL_47_DFFSR_184 gnd vdd FILL
XFILL_13_NAND3X1_127 gnd vdd FILL
XFILL_6_INVX1_7 gnd vdd FILL
XFILL_6_NOR2X1_169 gnd vdd FILL
XFILL_21_DFFSR_109 gnd vdd FILL
XFILL_12_NAND3X1_60 gnd vdd FILL
XFILL_47_DFFSR_195 gnd vdd FILL
XFILL_4_INVX1_30 gnd vdd FILL
XFILL_12_NAND3X1_71 gnd vdd FILL
XFILL_4_INVX1_41 gnd vdd FILL
XFILL_4_INVX1_52 gnd vdd FILL
XFILL_12_NAND3X1_82 gnd vdd FILL
XFILL_12_NAND3X1_93 gnd vdd FILL
XFILL_4_INVX1_63 gnd vdd FILL
XFILL_13_AOI22X1_2 gnd vdd FILL
XFILL_4_INVX1_74 gnd vdd FILL
XFILL_4_INVX1_85 gnd vdd FILL
XFILL_4_INVX1_96 gnd vdd FILL
XFILL_25_DFFSR_108 gnd vdd FILL
XFILL_25_DFFSR_119 gnd vdd FILL
XFILL_23_MUX2X1_105 gnd vdd FILL
XFILL_11_MUX2X1_6 gnd vdd FILL
XFILL_23_MUX2X1_116 gnd vdd FILL
XFILL_23_MUX2X1_127 gnd vdd FILL
XFILL_17_AOI22X1_1 gnd vdd FILL
XFILL_23_MUX2X1_138 gnd vdd FILL
XFILL_23_MUX2X1_149 gnd vdd FILL
XFILL_29_DFFSR_107 gnd vdd FILL
XFILL_6_MUX2X1_109 gnd vdd FILL
XFILL_19_DFFSR_10 gnd vdd FILL
XFILL_19_DFFSR_21 gnd vdd FILL
XFILL_2_BUFX4_50 gnd vdd FILL
XFILL_29_DFFSR_118 gnd vdd FILL
XFILL_2_BUFX4_61 gnd vdd FILL
XFILL_29_DFFSR_129 gnd vdd FILL
XFILL_19_DFFSR_32 gnd vdd FILL
XFILL_2_BUFX4_72 gnd vdd FILL
XFILL_2_BUFX4_83 gnd vdd FILL
XFILL_19_DFFSR_43 gnd vdd FILL
XFILL_3_OAI22X1_12 gnd vdd FILL
XFILL_19_DFFSR_54 gnd vdd FILL
XFILL_2_BUFX4_94 gnd vdd FILL
XFILL_19_DFFSR_65 gnd vdd FILL
XFILL_3_OAI22X1_23 gnd vdd FILL
XFILL_19_DFFSR_76 gnd vdd FILL
XFILL_3_OAI22X1_34 gnd vdd FILL
XFILL_19_DFFSR_87 gnd vdd FILL
XFILL_3_OAI22X1_45 gnd vdd FILL
XFILL_7_OAI21X1_14 gnd vdd FILL
XFILL_19_DFFSR_98 gnd vdd FILL
XFILL_7_OAI21X1_25 gnd vdd FILL
XFILL_59_DFFSR_20 gnd vdd FILL
XFILL_59_DFFSR_31 gnd vdd FILL
XFILL_59_DFFSR_42 gnd vdd FILL
XFILL_7_OAI21X1_36 gnd vdd FILL
XFILL_71_DFFSR_209 gnd vdd FILL
XFILL_7_OAI21X1_47 gnd vdd FILL
XFILL_59_DFFSR_53 gnd vdd FILL
XFILL_20_MUX2X1_4 gnd vdd FILL
XFILL_59_DFFSR_64 gnd vdd FILL
XFILL_59_DFFSR_75 gnd vdd FILL
XFILL_62_5_0 gnd vdd FILL
XFILL_59_DFFSR_86 gnd vdd FILL
XFILL_34_2_2 gnd vdd FILL
XFILL_25_NOR3X1_19 gnd vdd FILL
XFILL_59_DFFSR_97 gnd vdd FILL
XFILL_27_DFFSR_1 gnd vdd FILL
XFILL_75_DFFSR_208 gnd vdd FILL
XFILL_0_NOR2X1_203 gnd vdd FILL
XFILL_4_NOR2X1_7 gnd vdd FILL
XFILL_10_DFFSR_130 gnd vdd FILL
XFILL_75_DFFSR_219 gnd vdd FILL
XFILL_84_DFFSR_2 gnd vdd FILL
XFILL_10_DFFSR_141 gnd vdd FILL
XFILL_10_DFFSR_152 gnd vdd FILL
XFILL_6_NAND2X1_90 gnd vdd FILL
XFILL_28_DFFSR_30 gnd vdd FILL
XFILL_10_DFFSR_163 gnd vdd FILL
XFILL_10_DFFSR_174 gnd vdd FILL
XFILL_28_DFFSR_41 gnd vdd FILL
XFILL_29_NOR3X1_18 gnd vdd FILL
XFILL_12_2 gnd vdd FILL
XFILL_28_DFFSR_52 gnd vdd FILL
XFILL_10_DFFSR_185 gnd vdd FILL
XFILL_29_NOR3X1_29 gnd vdd FILL
XFILL_28_DFFSR_63 gnd vdd FILL
XFILL_14_CLKBUF1_10 gnd vdd FILL
XFILL_10_DFFSR_196 gnd vdd FILL
XFILL_14_CLKBUF1_21 gnd vdd FILL
XFILL_28_DFFSR_74 gnd vdd FILL
XFILL_79_DFFSR_207 gnd vdd FILL
XFILL_14_CLKBUF1_32 gnd vdd FILL
XFILL_28_DFFSR_85 gnd vdd FILL
XFILL_28_DFFSR_96 gnd vdd FILL
XFILL_79_DFFSR_218 gnd vdd FILL
XFILL_14_DFFSR_140 gnd vdd FILL
XFILL_79_DFFSR_229 gnd vdd FILL
XFILL_14_DFFSR_151 gnd vdd FILL
XFILL_14_DFFSR_162 gnd vdd FILL
XFILL_68_DFFSR_40 gnd vdd FILL
XFILL_14_DFFSR_173 gnd vdd FILL
XFILL_3_MUX2X1_5 gnd vdd FILL
XFILL_3_CLKBUF1_5 gnd vdd FILL
XFILL_68_DFFSR_51 gnd vdd FILL
XFILL_14_DFFSR_184 gnd vdd FILL
XFILL_68_DFFSR_62 gnd vdd FILL
XFILL_14_DFFSR_195 gnd vdd FILL
XFILL_68_DFFSR_73 gnd vdd FILL
XFILL_68_DFFSR_84 gnd vdd FILL
XFILL_11_DFFSR_7 gnd vdd FILL
XFILL_68_DFFSR_95 gnd vdd FILL
XFILL_18_DFFSR_150 gnd vdd FILL
XFILL_18_DFFSR_161 gnd vdd FILL
XFILL_18_DFFSR_172 gnd vdd FILL
XFILL_7_CLKBUF1_4 gnd vdd FILL
XFILL_49_DFFSR_5 gnd vdd FILL
XFILL_18_DFFSR_183 gnd vdd FILL
XFILL_18_DFFSR_194 gnd vdd FILL
XFILL_10_NOR3X1_30 gnd vdd FILL
XFILL_10_NOR3X1_41 gnd vdd FILL
XFILL_10_NOR3X1_52 gnd vdd FILL
XFILL_37_DFFSR_50 gnd vdd FILL
XFILL_37_DFFSR_61 gnd vdd FILL
XFILL_60_DFFSR_230 gnd vdd FILL
XFILL_37_DFFSR_72 gnd vdd FILL
XFILL_60_DFFSR_241 gnd vdd FILL
XFILL_37_DFFSR_83 gnd vdd FILL
XFILL_37_DFFSR_94 gnd vdd FILL
XFILL_60_DFFSR_252 gnd vdd FILL
XFILL_60_DFFSR_263 gnd vdd FILL
XFILL_60_DFFSR_274 gnd vdd FILL
XFILL_14_NOR3X1_40 gnd vdd FILL
XFILL_14_NOR3X1_51 gnd vdd FILL
XFILL_77_DFFSR_60 gnd vdd FILL
XFILL_77_DFFSR_71 gnd vdd FILL
XFILL_77_DFFSR_82 gnd vdd FILL
XFILL_64_DFFSR_240 gnd vdd FILL
XFILL_64_DFFSR_251 gnd vdd FILL
XFILL_77_DFFSR_93 gnd vdd FILL
XFILL_64_DFFSR_262 gnd vdd FILL
XFILL_64_DFFSR_273 gnd vdd FILL
XFILL_18_NOR3X1_50 gnd vdd FILL
XFILL_12_MUX2X1_101 gnd vdd FILL
XFILL_12_MUX2X1_112 gnd vdd FILL
XFILL_12_MUX2X1_123 gnd vdd FILL
XFILL_53_5_0 gnd vdd FILL
XFILL_0_2_2 gnd vdd FILL
XFILL_25_2_2 gnd vdd FILL
XFILL_12_MUX2X1_134 gnd vdd FILL
XFILL_17_NOR3X1_1 gnd vdd FILL
XFILL_12_MUX2X1_145 gnd vdd FILL
XFILL_68_DFFSR_250 gnd vdd FILL
XFILL_12_MUX2X1_156 gnd vdd FILL
XFILL_68_DFFSR_261 gnd vdd FILL
XFILL_12_MUX2X1_167 gnd vdd FILL
XFILL_23_CLKBUF1_2 gnd vdd FILL
XFILL_68_DFFSR_272 gnd vdd FILL
XFILL_12_MUX2X1_178 gnd vdd FILL
XFILL_46_DFFSR_70 gnd vdd FILL
XFILL_46_DFFSR_81 gnd vdd FILL
XFILL_46_DFFSR_92 gnd vdd FILL
XFILL_12_MUX2X1_189 gnd vdd FILL
XFILL_1_NOR2X1_12 gnd vdd FILL
XFILL_42_DFFSR_208 gnd vdd FILL
XFILL_1_NOR2X1_23 gnd vdd FILL
XFILL_42_DFFSR_219 gnd vdd FILL
XFILL_1_NOR2X1_34 gnd vdd FILL
XFILL_4_OAI21X1_9 gnd vdd FILL
XFILL_1_NOR2X1_45 gnd vdd FILL
XFILL_1_NOR2X1_56 gnd vdd FILL
XFILL_13_OAI21X1_50 gnd vdd FILL
XFILL_1_NOR2X1_67 gnd vdd FILL
XFILL_1_NOR2X1_78 gnd vdd FILL
XFILL_27_CLKBUF1_1 gnd vdd FILL
XFILL_86_DFFSR_80 gnd vdd FILL
XFILL_1_NOR2X1_89 gnd vdd FILL
XFILL_86_DFFSR_91 gnd vdd FILL
XFILL_5_NOR2X1_11 gnd vdd FILL
XFILL_46_DFFSR_207 gnd vdd FILL
XFILL_5_NOR2X1_22 gnd vdd FILL
XFILL_5_NOR2X1_33 gnd vdd FILL
XFILL_46_DFFSR_218 gnd vdd FILL
XFILL_8_OAI21X1_8 gnd vdd FILL
XFILL_46_DFFSR_229 gnd vdd FILL
XFILL_15_DFFSR_80 gnd vdd FILL
XFILL_5_NOR2X1_44 gnd vdd FILL
XFILL_5_NOR2X1_55 gnd vdd FILL
XFILL_15_DFFSR_91 gnd vdd FILL
XFILL_5_NOR2X1_66 gnd vdd FILL
XFILL_5_NOR2X1_77 gnd vdd FILL
XFILL_5_NOR2X1_88 gnd vdd FILL
XFILL_73_DFFSR_107 gnd vdd FILL
XFILL_5_NOR2X1_99 gnd vdd FILL
XFILL_9_NOR2X1_10 gnd vdd FILL
XFILL_73_DFFSR_118 gnd vdd FILL
XFILL_9_NOR2X1_21 gnd vdd FILL
XFILL_73_DFFSR_129 gnd vdd FILL
XFILL_9_NOR2X1_32 gnd vdd FILL
XFILL_9_NOR2X1_43 gnd vdd FILL
XFILL_55_DFFSR_90 gnd vdd FILL
XFILL_9_NOR2X1_54 gnd vdd FILL
XFILL_13_OAI22X1_5 gnd vdd FILL
XFILL_9_NOR2X1_65 gnd vdd FILL
XFILL_9_NOR2X1_76 gnd vdd FILL
XFILL_9_NOR2X1_87 gnd vdd FILL
XFILL_9_NOR2X1_98 gnd vdd FILL
XFILL_8_3_2 gnd vdd FILL
XFILL_77_DFFSR_106 gnd vdd FILL
XFILL_77_DFFSR_117 gnd vdd FILL
XFILL_2_MUX2X1_140 gnd vdd FILL
XFILL_77_DFFSR_128 gnd vdd FILL
XFILL_2_MUX2X1_151 gnd vdd FILL
XFILL_77_DFFSR_139 gnd vdd FILL
XFILL_2_MUX2X1_162 gnd vdd FILL
XFILL_17_OAI22X1_4 gnd vdd FILL
XFILL_15_NAND3X1_15 gnd vdd FILL
XFILL_2_MUX2X1_173 gnd vdd FILL
XFILL_15_NAND3X1_26 gnd vdd FILL
XFILL_15_NAND3X1_37 gnd vdd FILL
XFILL_2_MUX2X1_184 gnd vdd FILL
XFILL_15_NAND3X1_48 gnd vdd FILL
XFILL_15_NAND3X1_59 gnd vdd FILL
XFILL_35_CLKBUF1_15 gnd vdd FILL
XFILL_35_CLKBUF1_26 gnd vdd FILL
XFILL_35_CLKBUF1_37 gnd vdd FILL
XFILL_31_DFFSR_240 gnd vdd FILL
XFILL_31_DFFSR_251 gnd vdd FILL
XFILL_44_5_0 gnd vdd FILL
XFILL_31_DFFSR_262 gnd vdd FILL
XFILL_31_DFFSR_273 gnd vdd FILL
XFILL_16_2_2 gnd vdd FILL
XFILL_35_DFFSR_250 gnd vdd FILL
XFILL_11_BUFX4_18 gnd vdd FILL
XFILL_11_BUFX4_29 gnd vdd FILL
XFILL_35_DFFSR_261 gnd vdd FILL
XFILL_35_DFFSR_272 gnd vdd FILL
XFILL_1_MUX2X1_30 gnd vdd FILL
XFILL_7_DFFSR_90 gnd vdd FILL
XFILL_1_MUX2X1_41 gnd vdd FILL
XFILL_1_MUX2X1_52 gnd vdd FILL
XFILL_1_MUX2X1_63 gnd vdd FILL
XFILL_1_MUX2X1_74 gnd vdd FILL
XFILL_1_MUX2X1_85 gnd vdd FILL
XFILL_62_DFFSR_150 gnd vdd FILL
XFILL_62_DFFSR_161 gnd vdd FILL
XFILL_39_DFFSR_260 gnd vdd FILL
XFILL_14_NAND3X1_106 gnd vdd FILL
XFILL_1_MUX2X1_96 gnd vdd FILL
XFILL_62_DFFSR_172 gnd vdd FILL
XFILL_14_NAND3X1_117 gnd vdd FILL
XFILL_14_NAND3X1_128 gnd vdd FILL
XFILL_39_DFFSR_271 gnd vdd FILL
XFILL_62_DFFSR_183 gnd vdd FILL
XFILL_9_NAND2X1_9 gnd vdd FILL
XFILL_62_DFFSR_194 gnd vdd FILL
XFILL_5_MUX2X1_40 gnd vdd FILL
XFILL_13_DFFSR_207 gnd vdd FILL
XFILL_10_NAND3X1_7 gnd vdd FILL
XFILL_5_NAND3X1_10 gnd vdd FILL
XFILL_5_NAND3X1_21 gnd vdd FILL
XFILL_5_MUX2X1_51 gnd vdd FILL
XFILL_13_DFFSR_218 gnd vdd FILL
XFILL_5_MUX2X1_62 gnd vdd FILL
XFILL_13_DFFSR_229 gnd vdd FILL
XFILL_5_MUX2X1_73 gnd vdd FILL
XFILL_5_NAND3X1_32 gnd vdd FILL
XFILL_5_MUX2X1_84 gnd vdd FILL
XFILL_5_NAND3X1_43 gnd vdd FILL
XFILL_66_DFFSR_160 gnd vdd FILL
XFILL_5_MUX2X1_95 gnd vdd FILL
XFILL_5_NAND3X1_54 gnd vdd FILL
XFILL_50_DFFSR_5 gnd vdd FILL
XFILL_5_NAND3X1_65 gnd vdd FILL
XFILL_9_NAND2X1_12 gnd vdd FILL
XFILL_66_DFFSR_171 gnd vdd FILL
XFILL_9_NAND2X1_23 gnd vdd FILL
XFILL_5_NAND3X1_76 gnd vdd FILL
XFILL_66_DFFSR_182 gnd vdd FILL
XFILL_66_DFFSR_193 gnd vdd FILL
XFILL_9_NAND2X1_34 gnd vdd FILL
XFILL_40_DFFSR_107 gnd vdd FILL
XFILL_5_NAND3X1_87 gnd vdd FILL
XFILL_9_NAND2X1_45 gnd vdd FILL
XFILL_17_DFFSR_206 gnd vdd FILL
XFILL_40_DFFSR_118 gnd vdd FILL
XFILL_14_NAND3X1_6 gnd vdd FILL
XFILL_9_MUX2X1_50 gnd vdd FILL
XFILL_9_NAND2X1_56 gnd vdd FILL
XFILL_5_NAND3X1_98 gnd vdd FILL
XFILL_17_DFFSR_217 gnd vdd FILL
XFILL_17_DFFSR_228 gnd vdd FILL
XFILL_40_DFFSR_129 gnd vdd FILL
XFILL_9_MUX2X1_61 gnd vdd FILL
XFILL_9_NAND2X1_67 gnd vdd FILL
XFILL_9_NAND2X1_78 gnd vdd FILL
XFILL_5_INVX1_19 gnd vdd FILL
XFILL_17_DFFSR_239 gnd vdd FILL
XFILL_9_MUX2X1_72 gnd vdd FILL
XFILL_9_MUX2X1_83 gnd vdd FILL
XFILL_9_NAND2X1_89 gnd vdd FILL
XCLKBUF1_19 BUFX4_84/Y gnd DFFSR_84/CLK vdd CLKBUF1
XFILL_9_MUX2X1_94 gnd vdd FILL
XFILL_44_DFFSR_106 gnd vdd FILL
XFILL_67_3 gnd vdd FILL
XFILL_44_DFFSR_117 gnd vdd FILL
XFILL_44_DFFSR_128 gnd vdd FILL
XBUFX4_40 rst_n gnd BUFX4_54/A vdd BUFX4
XFILL_66_1_2 gnd vdd FILL
XBUFX4_51 rst_n gnd BUFX4_51/Y vdd BUFX4
XFILL_44_DFFSR_139 gnd vdd FILL
XFILL_12_AOI21X1_17 gnd vdd FILL
XBUFX4_62 rst_n gnd BUFX4_62/Y vdd BUFX4
XBUFX4_73 clk gnd BUFX4_73/Y vdd BUFX4
XFILL_12_AOI21X1_28 gnd vdd FILL
XBUFX4_84 clk gnd BUFX4_84/Y vdd BUFX4
XFILL_12_AOI21X1_39 gnd vdd FILL
XBUFX4_95 clk gnd BUFX4_95/Y vdd BUFX4
XFILL_48_DFFSR_105 gnd vdd FILL
XFILL_15_DFFSR_8 gnd vdd FILL
XFILL_48_DFFSR_116 gnd vdd FILL
XFILL_3_BUFX4_17 gnd vdd FILL
XFILL_48_DFFSR_127 gnd vdd FILL
XFILL_48_DFFSR_138 gnd vdd FILL
XFILL_3_BUFX4_28 gnd vdd FILL
XFILL_35_5_0 gnd vdd FILL
XFILL_72_DFFSR_9 gnd vdd FILL
XFILL_48_DFFSR_149 gnd vdd FILL
XFILL_3_BUFX4_39 gnd vdd FILL
XFILL_21_MUX2X1_60 gnd vdd FILL
XFILL_21_MUX2X1_71 gnd vdd FILL
XFILL_21_MUX2X1_82 gnd vdd FILL
XFILL_9_AOI22X1_10 gnd vdd FILL
XFILL_21_MUX2X1_93 gnd vdd FILL
XFILL_24_CLKBUF1_11 gnd vdd FILL
XFILL_24_CLKBUF1_22 gnd vdd FILL
XFILL_24_CLKBUF1_33 gnd vdd FILL
XFILL_0_NAND3X1_107 gnd vdd FILL
XFILL_0_NAND3X1_118 gnd vdd FILL
XFILL_0_NAND3X1_129 gnd vdd FILL
XFILL_7_CLKBUF1_15 gnd vdd FILL
XFILL_10_AND2X2_5 gnd vdd FILL
XFILL_7_CLKBUF1_26 gnd vdd FILL
XFILL_29_DFFSR_19 gnd vdd FILL
XFILL_7_CLKBUF1_37 gnd vdd FILL
XFILL_2_AOI21X1_12 gnd vdd FILL
XFILL_2_AOI21X1_23 gnd vdd FILL
XFILL_2_AOI21X1_34 gnd vdd FILL
XFILL_2_AOI21X1_45 gnd vdd FILL
XFILL_33_DFFSR_160 gnd vdd FILL
XFILL_12_OAI22X1_14 gnd vdd FILL
XFILL_2_AOI21X1_56 gnd vdd FILL
XFILL_33_DFFSR_171 gnd vdd FILL
XFILL_2_AOI21X1_67 gnd vdd FILL
XFILL_12_OAI22X1_25 gnd vdd FILL
XFILL_33_DFFSR_182 gnd vdd FILL
XFILL_2_AOI21X1_78 gnd vdd FILL
XFILL_33_DFFSR_193 gnd vdd FILL
XFILL_12_OAI22X1_36 gnd vdd FILL
XFILL_69_DFFSR_18 gnd vdd FILL
XFILL_12_OAI22X1_47 gnd vdd FILL
XFILL_69_DFFSR_29 gnd vdd FILL
XFILL_5_NOR2X1_100 gnd vdd FILL
XFILL_5_NOR2X1_111 gnd vdd FILL
XFILL_5_NOR2X1_122 gnd vdd FILL
XFILL_5_NOR2X1_133 gnd vdd FILL
XFILL_5_NOR2X1_144 gnd vdd FILL
XFILL_37_DFFSR_170 gnd vdd FILL
XFILL_5_NOR2X1_155 gnd vdd FILL
XFILL_5_NOR2X1_166 gnd vdd FILL
XFILL_37_DFFSR_181 gnd vdd FILL
XFILL_5_NOR2X1_177 gnd vdd FILL
XFILL_37_DFFSR_192 gnd vdd FILL
XFILL_11_DFFSR_106 gnd vdd FILL
XFILL_57_1_2 gnd vdd FILL
XFILL_5_NOR2X1_188 gnd vdd FILL
XFILL_11_DFFSR_117 gnd vdd FILL
XFILL_5_NOR2X1_199 gnd vdd FILL
XFILL_11_DFFSR_128 gnd vdd FILL
XFILL_11_NAND3X1_90 gnd vdd FILL
XFILL_11_DFFSR_139 gnd vdd FILL
XFILL_38_DFFSR_17 gnd vdd FILL
XFILL_38_DFFSR_28 gnd vdd FILL
XFILL_38_DFFSR_39 gnd vdd FILL
XFILL_26_5_0 gnd vdd FILL
XFILL_1_5_0 gnd vdd FILL
XFILL_15_DFFSR_105 gnd vdd FILL
XFILL_15_DFFSR_116 gnd vdd FILL
XFILL_22_MUX2X1_102 gnd vdd FILL
XFILL_15_DFFSR_127 gnd vdd FILL
XFILL_22_MUX2X1_113 gnd vdd FILL
XFILL_15_DFFSR_138 gnd vdd FILL
XFILL_22_MUX2X1_124 gnd vdd FILL
XFILL_78_DFFSR_16 gnd vdd FILL
XFILL_15_DFFSR_149 gnd vdd FILL
XFILL_22_MUX2X1_135 gnd vdd FILL
XFILL_10_AOI21X1_1 gnd vdd FILL
XFILL_78_DFFSR_27 gnd vdd FILL
XFILL_22_MUX2X1_146 gnd vdd FILL
XFILL_78_DFFSR_38 gnd vdd FILL
XFILL_78_DFFSR_49 gnd vdd FILL
XFILL_22_MUX2X1_157 gnd vdd FILL
XFILL_83_DFFSR_260 gnd vdd FILL
XFILL_22_MUX2X1_168 gnd vdd FILL
XFILL_19_DFFSR_104 gnd vdd FILL
XFILL_83_DFFSR_271 gnd vdd FILL
XFILL_40_0_2 gnd vdd FILL
XFILL_5_MUX2X1_106 gnd vdd FILL
XFILL_22_MUX2X1_179 gnd vdd FILL
XFILL_5_MUX2X1_117 gnd vdd FILL
XFILL_19_DFFSR_115 gnd vdd FILL
XFILL_19_DFFSR_126 gnd vdd FILL
XFILL_5_MUX2X1_128 gnd vdd FILL
XFILL_1_INVX1_12 gnd vdd FILL
XFILL_19_DFFSR_137 gnd vdd FILL
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
XFILL_5_MUX2X1_139 gnd vdd FILL
XFILL_1_INVX1_23 gnd vdd FILL
XFILL_1_INVX1_34 gnd vdd FILL
XFILL_19_DFFSR_148 gnd vdd FILL
XFILL_1_INVX1_45 gnd vdd FILL
XFILL_2_AND2X2_4 gnd vdd FILL
XFILL_1_INVX1_56 gnd vdd FILL
XFILL_2_OAI22X1_20 gnd vdd FILL
XFILL_19_DFFSR_159 gnd vdd FILL
XFILL_2_OAI22X1_31 gnd vdd FILL
XFILL_2_OAI22X1_42 gnd vdd FILL
XFILL_1_INVX1_67 gnd vdd FILL
XFILL_11_NOR3X1_17 gnd vdd FILL
XFILL_1_INVX1_78 gnd vdd FILL
XFILL_47_DFFSR_15 gnd vdd FILL
XFILL_6_OAI21X1_11 gnd vdd FILL
XFILL_87_DFFSR_270 gnd vdd FILL
XFILL_1_INVX1_89 gnd vdd FILL
XFILL_11_NOR3X1_28 gnd vdd FILL
XFILL_47_DFFSR_26 gnd vdd FILL
XFILL_11_NOR3X1_39 gnd vdd FILL
XFILL_6_OAI21X1_22 gnd vdd FILL
XFILL_47_DFFSR_37 gnd vdd FILL
XFILL_6_OAI21X1_33 gnd vdd FILL
XFILL_61_DFFSR_206 gnd vdd FILL
XFILL_47_DFFSR_48 gnd vdd FILL
XFILL_61_DFFSR_217 gnd vdd FILL
XFILL_6_OAI21X1_44 gnd vdd FILL
XFILL_47_DFFSR_59 gnd vdd FILL
XFILL_61_DFFSR_228 gnd vdd FILL
XFILL_61_DFFSR_239 gnd vdd FILL
XFILL_15_NOR3X1_16 gnd vdd FILL
XFILL_87_DFFSR_14 gnd vdd FILL
XFILL_15_NOR3X1_27 gnd vdd FILL
XFILL_87_DFFSR_25 gnd vdd FILL
XFILL_87_DFFSR_36 gnd vdd FILL
XFILL_15_NOR3X1_38 gnd vdd FILL
XFILL_32_DFFSR_2 gnd vdd FILL
XFILL_15_NOR3X1_49 gnd vdd FILL
XFILL_65_DFFSR_205 gnd vdd FILL
XFILL_87_DFFSR_47 gnd vdd FILL
XFILL_87_DFFSR_58 gnd vdd FILL
XFILL_65_DFFSR_216 gnd vdd FILL
XFILL_16_DFFSR_14 gnd vdd FILL
.ends

